library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.std_logic_unsigned.ALL;
entity street_image is
  port (clk_25   : in  std_logic;
        reset    : in  std_logic;
        vs_out   : out std_logic;
        hs_out   : out std_logic;
		  de_out   : out std_logic;
        r_out    : out std_logic_vector(1 downto 0);
        g_out    : out std_logic_vector(1 downto 0);
        b_out    : out std_logic_vector(1 downto 0));
end street_image;

architecture behave of street_image is

signal h_count   : std_logic_vector(9 downto 0) := "0000000000";
signal v_count   : std_logic_vector(9 downto 0) := "0000000000";
signal frame_num : std_logic_vector(9 downto 0) := "0000000000";
signal hs_1, vs_1, de_1 : std_logic;
signal new_frame : std_logic:='0';

type mem_typ is array(0 to 65535) of std_logic_vector(7 downto 0);
constant ROMINIT : mem_typ := (
0=>X"15",
1=>X"15",
2=>X"15",
3=>X"15",
4=>X"15",
5=>X"15",
6=>X"15",
7=>X"15",
8=>X"15",
9=>X"15",
10=>X"15",
11=>X"15",
12=>X"15",
13=>X"15",
14=>X"15",
15=>X"15",
16=>X"15",
17=>X"15",
18=>X"15",
19=>X"15",
20=>X"15",
21=>X"15",
22=>X"15",
23=>X"15",
24=>X"15",
25=>X"15",
26=>X"15",
27=>X"15",
28=>X"15",
29=>X"15",
30=>X"15",
31=>X"15",
32=>X"15",
33=>X"15",
34=>X"15",
35=>X"15",
36=>X"15",
37=>X"15",
38=>X"15",
39=>X"15",
40=>X"15",
41=>X"15",
42=>X"15",
43=>X"15",
44=>X"25",
45=>X"25",
46=>X"25",
47=>X"25",
48=>X"25",
49=>X"25",
50=>X"25",
51=>X"25",
52=>X"25",
53=>X"25",
54=>X"25",
55=>X"25",
56=>X"25",
57=>X"25",
58=>X"25",
59=>X"25",
60=>X"15",
61=>X"25",
62=>X"15",
63=>X"15",
64=>X"15",
65=>X"15",
66=>X"15",
67=>X"15",
68=>X"15",
69=>X"15",
70=>X"15",
71=>X"15",
72=>X"15",
73=>X"15",
74=>X"15",
75=>X"15",
76=>X"15",
77=>X"15",
78=>X"15",
79=>X"15",
80=>X"15",
81=>X"15",
82=>X"15",
83=>X"15",
84=>X"15",
85=>X"15",
86=>X"15",
87=>X"15",
88=>X"15",
89=>X"15",
90=>X"15",
91=>X"15",
92=>X"15",
93=>X"15",
94=>X"15",
95=>X"15",
96=>X"15",
97=>X"15",
98=>X"15",
99=>X"15",
100=>X"00",
101=>X"00",
102=>X"00",
103=>X"00",
104=>X"00",
105=>X"00",
106=>X"00",
107=>X"00",
108=>X"00",
109=>X"00",
110=>X"00",
111=>X"00",
112=>X"00",
113=>X"00",
114=>X"00",
115=>X"00",
116=>X"00",
117=>X"00",
118=>X"00",
119=>X"00",
120=>X"00",
121=>X"00",
122=>X"00",
123=>X"00",
124=>X"00",
125=>X"00",
126=>X"00",
127=>X"00",
128=>X"00",
129=>X"00",
130=>X"00",
131=>X"00",
132=>X"00",
133=>X"00",
134=>X"00",
135=>X"00",
136=>X"00",
137=>X"00",
138=>X"00",
139=>X"00",
140=>X"00",
141=>X"00",
142=>X"00",
143=>X"00",
144=>X"00",
145=>X"00",
146=>X"00",
147=>X"00",
148=>X"00",
149=>X"00",
150=>X"00",
151=>X"00",
152=>X"00",
153=>X"00",
154=>X"00",
155=>X"00",
156=>X"00",
157=>X"00",
158=>X"00",
159=>X"00",
160=>X"00",
161=>X"00",
162=>X"00",
163=>X"00",
164=>X"00",
165=>X"00",
166=>X"00",
167=>X"00",
168=>X"00",
169=>X"00",
170=>X"00",
171=>X"00",
172=>X"00",
173=>X"00",
174=>X"00",
175=>X"00",
176=>X"00",
177=>X"00",
178=>X"00",
179=>X"00",
180=>X"00",
181=>X"00",
182=>X"00",
183=>X"00",
184=>X"00",
185=>X"00",
186=>X"00",
187=>X"00",
188=>X"00",
189=>X"00",
190=>X"00",
191=>X"00",
192=>X"00",
193=>X"00",
194=>X"00",
195=>X"00",
196=>X"00",
197=>X"00",
198=>X"00",
199=>X"00",
200=>X"00",
201=>X"00",
202=>X"00",
203=>X"00",
204=>X"00",
205=>X"00",
206=>X"00",
207=>X"00",
208=>X"00",
209=>X"00",
210=>X"00",
211=>X"00",
212=>X"00",
213=>X"00",
214=>X"00",
215=>X"00",
216=>X"00",
217=>X"00",
218=>X"00",
219=>X"00",
220=>X"00",
221=>X"00",
222=>X"00",
223=>X"00",
224=>X"00",
225=>X"00",
226=>X"00",
227=>X"00",
228=>X"00",
229=>X"00",
230=>X"00",
231=>X"00",
232=>X"00",
233=>X"00",
234=>X"00",
235=>X"00",
236=>X"00",
237=>X"00",
238=>X"00",
239=>X"00",
240=>X"00",
241=>X"00",
242=>X"00",
243=>X"00",
244=>X"00",
245=>X"00",
246=>X"00",
247=>X"00",
248=>X"00",
249=>X"00",
250=>X"00",
251=>X"00",
252=>X"00",
253=>X"00",
254=>X"00",
255=>X"00",
256=>X"15",
257=>X"15",
258=>X"15",
259=>X"15",
260=>X"15",
261=>X"15",
262=>X"15",
263=>X"15",
264=>X"15",
265=>X"15",
266=>X"15",
267=>X"15",
268=>X"15",
269=>X"15",
270=>X"15",
271=>X"15",
272=>X"15",
273=>X"15",
274=>X"15",
275=>X"15",
276=>X"15",
277=>X"15",
278=>X"15",
279=>X"15",
280=>X"15",
281=>X"15",
282=>X"15",
283=>X"15",
284=>X"15",
285=>X"15",
286=>X"15",
287=>X"15",
288=>X"15",
289=>X"15",
290=>X"15",
291=>X"15",
292=>X"15",
293=>X"15",
294=>X"15",
295=>X"15",
296=>X"25",
297=>X"15",
298=>X"25",
299=>X"15",
300=>X"25",
301=>X"25",
302=>X"25",
303=>X"25",
304=>X"25",
305=>X"25",
306=>X"25",
307=>X"25",
308=>X"25",
309=>X"25",
310=>X"25",
311=>X"25",
312=>X"25",
313=>X"25",
314=>X"25",
315=>X"25",
316=>X"25",
317=>X"15",
318=>X"25",
319=>X"15",
320=>X"25",
321=>X"15",
322=>X"15",
323=>X"15",
324=>X"15",
325=>X"15",
326=>X"15",
327=>X"15",
328=>X"15",
329=>X"15",
330=>X"15",
331=>X"15",
332=>X"15",
333=>X"15",
334=>X"15",
335=>X"15",
336=>X"15",
337=>X"15",
338=>X"15",
339=>X"15",
340=>X"15",
341=>X"15",
342=>X"15",
343=>X"15",
344=>X"15",
345=>X"15",
346=>X"15",
347=>X"15",
348=>X"15",
349=>X"15",
350=>X"15",
351=>X"15",
352=>X"15",
353=>X"15",
354=>X"15",
355=>X"15",
356=>X"00",
357=>X"00",
358=>X"00",
359=>X"00",
360=>X"00",
361=>X"00",
362=>X"00",
363=>X"00",
364=>X"00",
365=>X"00",
366=>X"00",
367=>X"00",
368=>X"00",
369=>X"00",
370=>X"00",
371=>X"00",
372=>X"00",
373=>X"00",
374=>X"00",
375=>X"00",
376=>X"00",
377=>X"00",
378=>X"00",
379=>X"00",
380=>X"00",
381=>X"00",
382=>X"00",
383=>X"00",
384=>X"00",
385=>X"00",
386=>X"00",
387=>X"00",
388=>X"00",
389=>X"00",
390=>X"00",
391=>X"00",
392=>X"00",
393=>X"00",
394=>X"00",
395=>X"00",
396=>X"00",
397=>X"00",
398=>X"00",
399=>X"00",
400=>X"00",
401=>X"00",
402=>X"00",
403=>X"00",
404=>X"00",
405=>X"00",
406=>X"00",
407=>X"00",
408=>X"00",
409=>X"00",
410=>X"00",
411=>X"00",
412=>X"00",
413=>X"00",
414=>X"00",
415=>X"00",
416=>X"00",
417=>X"00",
418=>X"00",
419=>X"00",
420=>X"00",
421=>X"00",
422=>X"00",
423=>X"00",
424=>X"00",
425=>X"00",
426=>X"00",
427=>X"00",
428=>X"00",
429=>X"00",
430=>X"00",
431=>X"00",
432=>X"00",
433=>X"00",
434=>X"00",
435=>X"00",
436=>X"00",
437=>X"00",
438=>X"00",
439=>X"00",
440=>X"00",
441=>X"00",
442=>X"00",
443=>X"00",
444=>X"00",
445=>X"00",
446=>X"00",
447=>X"00",
448=>X"00",
449=>X"00",
450=>X"00",
451=>X"00",
452=>X"00",
453=>X"00",
454=>X"00",
455=>X"00",
456=>X"00",
457=>X"00",
458=>X"00",
459=>X"00",
460=>X"00",
461=>X"00",
462=>X"00",
463=>X"00",
464=>X"00",
465=>X"00",
466=>X"00",
467=>X"00",
468=>X"00",
469=>X"00",
470=>X"00",
471=>X"00",
472=>X"00",
473=>X"00",
474=>X"00",
475=>X"00",
476=>X"00",
477=>X"00",
478=>X"00",
479=>X"00",
480=>X"00",
481=>X"00",
482=>X"00",
483=>X"00",
484=>X"00",
485=>X"00",
486=>X"00",
487=>X"00",
488=>X"00",
489=>X"00",
490=>X"00",
491=>X"00",
492=>X"00",
493=>X"00",
494=>X"00",
495=>X"00",
496=>X"00",
497=>X"00",
498=>X"00",
499=>X"00",
500=>X"00",
501=>X"00",
502=>X"00",
503=>X"00",
504=>X"00",
505=>X"00",
506=>X"00",
507=>X"00",
508=>X"00",
509=>X"00",
510=>X"00",
511=>X"00",
512=>X"15",
513=>X"15",
514=>X"15",
515=>X"15",
516=>X"15",
517=>X"15",
518=>X"15",
519=>X"15",
520=>X"15",
521=>X"15",
522=>X"15",
523=>X"15",
524=>X"15",
525=>X"15",
526=>X"15",
527=>X"15",
528=>X"15",
529=>X"15",
530=>X"15",
531=>X"15",
532=>X"15",
533=>X"15",
534=>X"15",
535=>X"15",
536=>X"15",
537=>X"15",
538=>X"15",
539=>X"15",
540=>X"15",
541=>X"15",
542=>X"15",
543=>X"15",
544=>X"15",
545=>X"15",
546=>X"15",
547=>X"15",
548=>X"15",
549=>X"15",
550=>X"15",
551=>X"15",
552=>X"15",
553=>X"15",
554=>X"15",
555=>X"15",
556=>X"15",
557=>X"15",
558=>X"25",
559=>X"25",
560=>X"25",
561=>X"25",
562=>X"25",
563=>X"25",
564=>X"25",
565=>X"25",
566=>X"25",
567=>X"25",
568=>X"25",
569=>X"25",
570=>X"25",
571=>X"25",
572=>X"25",
573=>X"25",
574=>X"15",
575=>X"15",
576=>X"15",
577=>X"15",
578=>X"15",
579=>X"15",
580=>X"15",
581=>X"15",
582=>X"15",
583=>X"15",
584=>X"15",
585=>X"15",
586=>X"15",
587=>X"15",
588=>X"15",
589=>X"15",
590=>X"15",
591=>X"15",
592=>X"15",
593=>X"15",
594=>X"15",
595=>X"15",
596=>X"15",
597=>X"15",
598=>X"15",
599=>X"15",
600=>X"15",
601=>X"15",
602=>X"15",
603=>X"15",
604=>X"15",
605=>X"15",
606=>X"15",
607=>X"15",
608=>X"15",
609=>X"15",
610=>X"15",
611=>X"15",
612=>X"00",
613=>X"00",
614=>X"00",
615=>X"00",
616=>X"00",
617=>X"00",
618=>X"00",
619=>X"00",
620=>X"00",
621=>X"00",
622=>X"00",
623=>X"00",
624=>X"00",
625=>X"00",
626=>X"00",
627=>X"00",
628=>X"00",
629=>X"00",
630=>X"00",
631=>X"00",
632=>X"00",
633=>X"00",
634=>X"00",
635=>X"00",
636=>X"00",
637=>X"00",
638=>X"00",
639=>X"00",
640=>X"00",
641=>X"00",
642=>X"00",
643=>X"00",
644=>X"00",
645=>X"00",
646=>X"00",
647=>X"00",
648=>X"00",
649=>X"00",
650=>X"00",
651=>X"00",
652=>X"00",
653=>X"00",
654=>X"00",
655=>X"00",
656=>X"00",
657=>X"00",
658=>X"00",
659=>X"00",
660=>X"00",
661=>X"00",
662=>X"00",
663=>X"00",
664=>X"00",
665=>X"00",
666=>X"00",
667=>X"00",
668=>X"00",
669=>X"00",
670=>X"00",
671=>X"00",
672=>X"00",
673=>X"00",
674=>X"00",
675=>X"00",
676=>X"00",
677=>X"00",
678=>X"00",
679=>X"00",
680=>X"00",
681=>X"00",
682=>X"00",
683=>X"00",
684=>X"00",
685=>X"00",
686=>X"00",
687=>X"00",
688=>X"00",
689=>X"00",
690=>X"00",
691=>X"00",
692=>X"00",
693=>X"00",
694=>X"00",
695=>X"00",
696=>X"00",
697=>X"00",
698=>X"00",
699=>X"00",
700=>X"00",
701=>X"00",
702=>X"00",
703=>X"00",
704=>X"00",
705=>X"00",
706=>X"00",
707=>X"00",
708=>X"00",
709=>X"00",
710=>X"00",
711=>X"00",
712=>X"00",
713=>X"00",
714=>X"00",
715=>X"00",
716=>X"00",
717=>X"00",
718=>X"00",
719=>X"00",
720=>X"00",
721=>X"00",
722=>X"00",
723=>X"00",
724=>X"00",
725=>X"00",
726=>X"00",
727=>X"00",
728=>X"00",
729=>X"00",
730=>X"00",
731=>X"00",
732=>X"00",
733=>X"00",
734=>X"00",
735=>X"00",
736=>X"00",
737=>X"00",
738=>X"00",
739=>X"00",
740=>X"00",
741=>X"00",
742=>X"00",
743=>X"00",
744=>X"00",
745=>X"00",
746=>X"00",
747=>X"00",
748=>X"00",
749=>X"00",
750=>X"00",
751=>X"00",
752=>X"00",
753=>X"00",
754=>X"00",
755=>X"00",
756=>X"00",
757=>X"00",
758=>X"00",
759=>X"00",
760=>X"00",
761=>X"00",
762=>X"00",
763=>X"00",
764=>X"00",
765=>X"00",
766=>X"00",
767=>X"00",
768=>X"15",
769=>X"15",
770=>X"15",
771=>X"15",
772=>X"15",
773=>X"15",
774=>X"15",
775=>X"15",
776=>X"15",
777=>X"15",
778=>X"15",
779=>X"15",
780=>X"15",
781=>X"15",
782=>X"15",
783=>X"15",
784=>X"15",
785=>X"15",
786=>X"15",
787=>X"15",
788=>X"15",
789=>X"15",
790=>X"15",
791=>X"15",
792=>X"15",
793=>X"15",
794=>X"15",
795=>X"15",
796=>X"15",
797=>X"15",
798=>X"15",
799=>X"15",
800=>X"15",
801=>X"15",
802=>X"15",
803=>X"15",
804=>X"15",
805=>X"15",
806=>X"15",
807=>X"15",
808=>X"15",
809=>X"15",
810=>X"25",
811=>X"15",
812=>X"15",
813=>X"25",
814=>X"25",
815=>X"25",
816=>X"25",
817=>X"25",
818=>X"25",
819=>X"25",
820=>X"25",
821=>X"25",
822=>X"25",
823=>X"25",
824=>X"25",
825=>X"25",
826=>X"25",
827=>X"15",
828=>X"25",
829=>X"25",
830=>X"25",
831=>X"15",
832=>X"25",
833=>X"15",
834=>X"15",
835=>X"15",
836=>X"15",
837=>X"15",
838=>X"15",
839=>X"15",
840=>X"15",
841=>X"15",
842=>X"15",
843=>X"15",
844=>X"15",
845=>X"15",
846=>X"15",
847=>X"15",
848=>X"15",
849=>X"15",
850=>X"15",
851=>X"15",
852=>X"15",
853=>X"15",
854=>X"15",
855=>X"15",
856=>X"15",
857=>X"15",
858=>X"15",
859=>X"15",
860=>X"15",
861=>X"15",
862=>X"15",
863=>X"15",
864=>X"15",
865=>X"15",
866=>X"15",
867=>X"15",
868=>X"00",
869=>X"00",
870=>X"00",
871=>X"00",
872=>X"00",
873=>X"00",
874=>X"00",
875=>X"00",
876=>X"00",
877=>X"00",
878=>X"00",
879=>X"00",
880=>X"00",
881=>X"00",
882=>X"00",
883=>X"00",
884=>X"00",
885=>X"00",
886=>X"00",
887=>X"00",
888=>X"00",
889=>X"00",
890=>X"00",
891=>X"00",
892=>X"00",
893=>X"00",
894=>X"00",
895=>X"00",
896=>X"00",
897=>X"00",
898=>X"00",
899=>X"00",
900=>X"00",
901=>X"00",
902=>X"00",
903=>X"00",
904=>X"00",
905=>X"00",
906=>X"00",
907=>X"00",
908=>X"00",
909=>X"00",
910=>X"00",
911=>X"00",
912=>X"00",
913=>X"00",
914=>X"00",
915=>X"00",
916=>X"00",
917=>X"00",
918=>X"00",
919=>X"00",
920=>X"00",
921=>X"00",
922=>X"00",
923=>X"00",
924=>X"00",
925=>X"00",
926=>X"00",
927=>X"00",
928=>X"00",
929=>X"00",
930=>X"00",
931=>X"00",
932=>X"00",
933=>X"00",
934=>X"00",
935=>X"00",
936=>X"00",
937=>X"00",
938=>X"00",
939=>X"00",
940=>X"00",
941=>X"00",
942=>X"00",
943=>X"00",
944=>X"00",
945=>X"00",
946=>X"00",
947=>X"00",
948=>X"00",
949=>X"00",
950=>X"00",
951=>X"00",
952=>X"00",
953=>X"00",
954=>X"00",
955=>X"00",
956=>X"00",
957=>X"00",
958=>X"00",
959=>X"00",
960=>X"00",
961=>X"00",
962=>X"00",
963=>X"00",
964=>X"00",
965=>X"00",
966=>X"00",
967=>X"00",
968=>X"00",
969=>X"00",
970=>X"00",
971=>X"00",
972=>X"00",
973=>X"00",
974=>X"00",
975=>X"00",
976=>X"00",
977=>X"00",
978=>X"00",
979=>X"00",
980=>X"00",
981=>X"00",
982=>X"00",
983=>X"00",
984=>X"00",
985=>X"00",
986=>X"00",
987=>X"00",
988=>X"00",
989=>X"00",
990=>X"00",
991=>X"00",
992=>X"00",
993=>X"00",
994=>X"00",
995=>X"00",
996=>X"00",
997=>X"00",
998=>X"00",
999=>X"00",
1000=>X"00",
1001=>X"00",
1002=>X"00",
1003=>X"00",
1004=>X"00",
1005=>X"00",
1006=>X"00",
1007=>X"00",
1008=>X"00",
1009=>X"00",
1010=>X"00",
1011=>X"00",
1012=>X"00",
1013=>X"00",
1014=>X"00",
1015=>X"00",
1016=>X"00",
1017=>X"00",
1018=>X"00",
1019=>X"00",
1020=>X"00",
1021=>X"00",
1022=>X"00",
1023=>X"00",
1024=>X"15",
1025=>X"15",
1026=>X"15",
1027=>X"15",
1028=>X"15",
1029=>X"15",
1030=>X"15",
1031=>X"15",
1032=>X"15",
1033=>X"15",
1034=>X"15",
1035=>X"15",
1036=>X"15",
1037=>X"15",
1038=>X"15",
1039=>X"15",
1040=>X"15",
1041=>X"15",
1042=>X"15",
1043=>X"15",
1044=>X"15",
1045=>X"15",
1046=>X"15",
1047=>X"15",
1048=>X"15",
1049=>X"15",
1050=>X"15",
1051=>X"15",
1052=>X"15",
1053=>X"15",
1054=>X"15",
1055=>X"15",
1056=>X"15",
1057=>X"15",
1058=>X"15",
1059=>X"15",
1060=>X"15",
1061=>X"15",
1062=>X"15",
1063=>X"15",
1064=>X"25",
1065=>X"15",
1066=>X"15",
1067=>X"15",
1068=>X"25",
1069=>X"25",
1070=>X"25",
1071=>X"25",
1072=>X"25",
1073=>X"25",
1074=>X"25",
1075=>X"25",
1076=>X"25",
1077=>X"25",
1078=>X"25",
1079=>X"25",
1080=>X"25",
1081=>X"25",
1082=>X"25",
1083=>X"15",
1084=>X"15",
1085=>X"15",
1086=>X"15",
1087=>X"15",
1088=>X"15",
1089=>X"15",
1090=>X"25",
1091=>X"15",
1092=>X"15",
1093=>X"15",
1094=>X"15",
1095=>X"15",
1096=>X"15",
1097=>X"15",
1098=>X"15",
1099=>X"15",
1100=>X"15",
1101=>X"15",
1102=>X"15",
1103=>X"15",
1104=>X"15",
1105=>X"15",
1106=>X"15",
1107=>X"15",
1108=>X"15",
1109=>X"15",
1110=>X"15",
1111=>X"15",
1112=>X"15",
1113=>X"15",
1114=>X"15",
1115=>X"15",
1116=>X"15",
1117=>X"15",
1118=>X"15",
1119=>X"15",
1120=>X"15",
1121=>X"15",
1122=>X"15",
1123=>X"15",
1124=>X"00",
1125=>X"00",
1126=>X"00",
1127=>X"00",
1128=>X"00",
1129=>X"00",
1130=>X"00",
1131=>X"00",
1132=>X"00",
1133=>X"00",
1134=>X"00",
1135=>X"00",
1136=>X"00",
1137=>X"00",
1138=>X"00",
1139=>X"00",
1140=>X"00",
1141=>X"00",
1142=>X"00",
1143=>X"00",
1144=>X"00",
1145=>X"00",
1146=>X"00",
1147=>X"00",
1148=>X"00",
1149=>X"00",
1150=>X"00",
1151=>X"00",
1152=>X"00",
1153=>X"00",
1154=>X"00",
1155=>X"00",
1156=>X"00",
1157=>X"00",
1158=>X"00",
1159=>X"00",
1160=>X"00",
1161=>X"00",
1162=>X"00",
1163=>X"00",
1164=>X"00",
1165=>X"00",
1166=>X"00",
1167=>X"00",
1168=>X"00",
1169=>X"00",
1170=>X"00",
1171=>X"00",
1172=>X"00",
1173=>X"00",
1174=>X"00",
1175=>X"00",
1176=>X"00",
1177=>X"00",
1178=>X"00",
1179=>X"00",
1180=>X"00",
1181=>X"00",
1182=>X"00",
1183=>X"00",
1184=>X"00",
1185=>X"00",
1186=>X"00",
1187=>X"00",
1188=>X"00",
1189=>X"00",
1190=>X"00",
1191=>X"00",
1192=>X"00",
1193=>X"00",
1194=>X"00",
1195=>X"00",
1196=>X"00",
1197=>X"00",
1198=>X"00",
1199=>X"00",
1200=>X"00",
1201=>X"00",
1202=>X"00",
1203=>X"00",
1204=>X"00",
1205=>X"00",
1206=>X"00",
1207=>X"00",
1208=>X"00",
1209=>X"00",
1210=>X"00",
1211=>X"00",
1212=>X"00",
1213=>X"00",
1214=>X"00",
1215=>X"00",
1216=>X"00",
1217=>X"00",
1218=>X"00",
1219=>X"00",
1220=>X"00",
1221=>X"00",
1222=>X"00",
1223=>X"00",
1224=>X"00",
1225=>X"00",
1226=>X"00",
1227=>X"00",
1228=>X"00",
1229=>X"00",
1230=>X"00",
1231=>X"00",
1232=>X"00",
1233=>X"00",
1234=>X"00",
1235=>X"00",
1236=>X"00",
1237=>X"00",
1238=>X"00",
1239=>X"00",
1240=>X"00",
1241=>X"00",
1242=>X"00",
1243=>X"00",
1244=>X"00",
1245=>X"00",
1246=>X"00",
1247=>X"00",
1248=>X"00",
1249=>X"00",
1250=>X"00",
1251=>X"00",
1252=>X"00",
1253=>X"00",
1254=>X"00",
1255=>X"00",
1256=>X"00",
1257=>X"00",
1258=>X"00",
1259=>X"00",
1260=>X"00",
1261=>X"00",
1262=>X"00",
1263=>X"00",
1264=>X"00",
1265=>X"00",
1266=>X"00",
1267=>X"00",
1268=>X"00",
1269=>X"00",
1270=>X"00",
1271=>X"00",
1272=>X"00",
1273=>X"00",
1274=>X"00",
1275=>X"00",
1276=>X"00",
1277=>X"00",
1278=>X"00",
1279=>X"00",
1280=>X"15",
1281=>X"15",
1282=>X"15",
1283=>X"15",
1284=>X"15",
1285=>X"15",
1286=>X"15",
1287=>X"15",
1288=>X"15",
1289=>X"15",
1290=>X"15",
1291=>X"15",
1292=>X"15",
1293=>X"15",
1294=>X"15",
1295=>X"15",
1296=>X"15",
1297=>X"15",
1298=>X"15",
1299=>X"15",
1300=>X"15",
1301=>X"15",
1302=>X"15",
1303=>X"15",
1304=>X"15",
1305=>X"15",
1306=>X"15",
1307=>X"15",
1308=>X"15",
1309=>X"15",
1310=>X"15",
1311=>X"15",
1312=>X"15",
1313=>X"15",
1314=>X"15",
1315=>X"15",
1316=>X"15",
1317=>X"15",
1318=>X"15",
1319=>X"15",
1320=>X"25",
1321=>X"15",
1322=>X"15",
1323=>X"15",
1324=>X"25",
1325=>X"25",
1326=>X"25",
1327=>X"25",
1328=>X"25",
1329=>X"25",
1330=>X"25",
1331=>X"25",
1332=>X"25",
1333=>X"25",
1334=>X"25",
1335=>X"25",
1336=>X"25",
1337=>X"25",
1338=>X"25",
1339=>X"25",
1340=>X"25",
1341=>X"25",
1342=>X"25",
1343=>X"25",
1344=>X"25",
1345=>X"15",
1346=>X"25",
1347=>X"15",
1348=>X"25",
1349=>X"15",
1350=>X"15",
1351=>X"25",
1352=>X"15",
1353=>X"15",
1354=>X"15",
1355=>X"15",
1356=>X"15",
1357=>X"15",
1358=>X"15",
1359=>X"15",
1360=>X"15",
1361=>X"15",
1362=>X"15",
1363=>X"15",
1364=>X"15",
1365=>X"15",
1366=>X"15",
1367=>X"15",
1368=>X"15",
1369=>X"15",
1370=>X"15",
1371=>X"15",
1372=>X"15",
1373=>X"15",
1374=>X"15",
1375=>X"15",
1376=>X"15",
1377=>X"15",
1378=>X"15",
1379=>X"15",
1380=>X"00",
1381=>X"00",
1382=>X"00",
1383=>X"00",
1384=>X"00",
1385=>X"00",
1386=>X"00",
1387=>X"00",
1388=>X"00",
1389=>X"00",
1390=>X"00",
1391=>X"00",
1392=>X"00",
1393=>X"00",
1394=>X"00",
1395=>X"00",
1396=>X"00",
1397=>X"00",
1398=>X"00",
1399=>X"00",
1400=>X"00",
1401=>X"00",
1402=>X"00",
1403=>X"00",
1404=>X"00",
1405=>X"00",
1406=>X"00",
1407=>X"00",
1408=>X"00",
1409=>X"00",
1410=>X"00",
1411=>X"00",
1412=>X"00",
1413=>X"00",
1414=>X"00",
1415=>X"00",
1416=>X"00",
1417=>X"00",
1418=>X"00",
1419=>X"00",
1420=>X"00",
1421=>X"00",
1422=>X"00",
1423=>X"00",
1424=>X"00",
1425=>X"00",
1426=>X"00",
1427=>X"00",
1428=>X"00",
1429=>X"00",
1430=>X"00",
1431=>X"00",
1432=>X"00",
1433=>X"00",
1434=>X"00",
1435=>X"00",
1436=>X"00",
1437=>X"00",
1438=>X"00",
1439=>X"00",
1440=>X"00",
1441=>X"00",
1442=>X"00",
1443=>X"00",
1444=>X"00",
1445=>X"00",
1446=>X"00",
1447=>X"00",
1448=>X"00",
1449=>X"00",
1450=>X"00",
1451=>X"00",
1452=>X"00",
1453=>X"00",
1454=>X"00",
1455=>X"00",
1456=>X"00",
1457=>X"00",
1458=>X"00",
1459=>X"00",
1460=>X"00",
1461=>X"00",
1462=>X"00",
1463=>X"00",
1464=>X"00",
1465=>X"00",
1466=>X"00",
1467=>X"00",
1468=>X"00",
1469=>X"00",
1470=>X"00",
1471=>X"00",
1472=>X"00",
1473=>X"00",
1474=>X"00",
1475=>X"00",
1476=>X"00",
1477=>X"00",
1478=>X"00",
1479=>X"00",
1480=>X"00",
1481=>X"00",
1482=>X"00",
1483=>X"00",
1484=>X"00",
1485=>X"00",
1486=>X"00",
1487=>X"00",
1488=>X"00",
1489=>X"00",
1490=>X"00",
1491=>X"00",
1492=>X"00",
1493=>X"00",
1494=>X"00",
1495=>X"00",
1496=>X"00",
1497=>X"00",
1498=>X"00",
1499=>X"00",
1500=>X"00",
1501=>X"00",
1502=>X"00",
1503=>X"00",
1504=>X"00",
1505=>X"00",
1506=>X"00",
1507=>X"00",
1508=>X"00",
1509=>X"00",
1510=>X"00",
1511=>X"00",
1512=>X"00",
1513=>X"00",
1514=>X"00",
1515=>X"00",
1516=>X"00",
1517=>X"00",
1518=>X"00",
1519=>X"00",
1520=>X"00",
1521=>X"00",
1522=>X"00",
1523=>X"00",
1524=>X"00",
1525=>X"00",
1526=>X"00",
1527=>X"00",
1528=>X"00",
1529=>X"00",
1530=>X"00",
1531=>X"00",
1532=>X"00",
1533=>X"00",
1534=>X"00",
1535=>X"00",
1536=>X"15",
1537=>X"15",
1538=>X"15",
1539=>X"15",
1540=>X"15",
1541=>X"15",
1542=>X"15",
1543=>X"15",
1544=>X"15",
1545=>X"15",
1546=>X"15",
1547=>X"15",
1548=>X"15",
1549=>X"15",
1550=>X"15",
1551=>X"15",
1552=>X"15",
1553=>X"15",
1554=>X"15",
1555=>X"15",
1556=>X"15",
1557=>X"15",
1558=>X"15",
1559=>X"15",
1560=>X"15",
1561=>X"15",
1562=>X"15",
1563=>X"15",
1564=>X"15",
1565=>X"15",
1566=>X"15",
1567=>X"15",
1568=>X"15",
1569=>X"15",
1570=>X"15",
1571=>X"15",
1572=>X"15",
1573=>X"15",
1574=>X"15",
1575=>X"15",
1576=>X"25",
1577=>X"15",
1578=>X"25",
1579=>X"15",
1580=>X"25",
1581=>X"25",
1582=>X"25",
1583=>X"25",
1584=>X"25",
1585=>X"25",
1586=>X"25",
1587=>X"25",
1588=>X"25",
1589=>X"25",
1590=>X"25",
1591=>X"25",
1592=>X"25",
1593=>X"25",
1594=>X"25",
1595=>X"25",
1596=>X"25",
1597=>X"25",
1598=>X"25",
1599=>X"25",
1600=>X"25",
1601=>X"15",
1602=>X"15",
1603=>X"15",
1604=>X"25",
1605=>X"25",
1606=>X"15",
1607=>X"25",
1608=>X"15",
1609=>X"25",
1610=>X"15",
1611=>X"15",
1612=>X"25",
1613=>X"15",
1614=>X"15",
1615=>X"15",
1616=>X"15",
1617=>X"15",
1618=>X"15",
1619=>X"15",
1620=>X"15",
1621=>X"15",
1622=>X"15",
1623=>X"15",
1624=>X"15",
1625=>X"15",
1626=>X"15",
1627=>X"15",
1628=>X"15",
1629=>X"15",
1630=>X"15",
1631=>X"15",
1632=>X"15",
1633=>X"15",
1634=>X"15",
1635=>X"15",
1636=>X"00",
1637=>X"00",
1638=>X"00",
1639=>X"00",
1640=>X"00",
1641=>X"00",
1642=>X"00",
1643=>X"00",
1644=>X"00",
1645=>X"00",
1646=>X"00",
1647=>X"00",
1648=>X"00",
1649=>X"00",
1650=>X"00",
1651=>X"00",
1652=>X"00",
1653=>X"00",
1654=>X"00",
1655=>X"00",
1656=>X"00",
1657=>X"00",
1658=>X"00",
1659=>X"00",
1660=>X"00",
1661=>X"00",
1662=>X"00",
1663=>X"00",
1664=>X"00",
1665=>X"00",
1666=>X"00",
1667=>X"00",
1668=>X"00",
1669=>X"00",
1670=>X"00",
1671=>X"00",
1672=>X"00",
1673=>X"00",
1674=>X"00",
1675=>X"00",
1676=>X"00",
1677=>X"00",
1678=>X"00",
1679=>X"00",
1680=>X"00",
1681=>X"00",
1682=>X"00",
1683=>X"00",
1684=>X"00",
1685=>X"00",
1686=>X"00",
1687=>X"00",
1688=>X"00",
1689=>X"00",
1690=>X"00",
1691=>X"00",
1692=>X"00",
1693=>X"00",
1694=>X"00",
1695=>X"00",
1696=>X"00",
1697=>X"00",
1698=>X"00",
1699=>X"00",
1700=>X"00",
1701=>X"00",
1702=>X"00",
1703=>X"00",
1704=>X"00",
1705=>X"00",
1706=>X"00",
1707=>X"00",
1708=>X"00",
1709=>X"00",
1710=>X"00",
1711=>X"00",
1712=>X"00",
1713=>X"00",
1714=>X"00",
1715=>X"00",
1716=>X"00",
1717=>X"00",
1718=>X"00",
1719=>X"00",
1720=>X"00",
1721=>X"00",
1722=>X"00",
1723=>X"00",
1724=>X"00",
1725=>X"00",
1726=>X"00",
1727=>X"00",
1728=>X"00",
1729=>X"00",
1730=>X"00",
1731=>X"00",
1732=>X"00",
1733=>X"00",
1734=>X"00",
1735=>X"00",
1736=>X"00",
1737=>X"00",
1738=>X"00",
1739=>X"00",
1740=>X"00",
1741=>X"00",
1742=>X"00",
1743=>X"00",
1744=>X"00",
1745=>X"00",
1746=>X"00",
1747=>X"00",
1748=>X"00",
1749=>X"00",
1750=>X"00",
1751=>X"00",
1752=>X"00",
1753=>X"00",
1754=>X"00",
1755=>X"00",
1756=>X"00",
1757=>X"00",
1758=>X"00",
1759=>X"00",
1760=>X"00",
1761=>X"00",
1762=>X"00",
1763=>X"00",
1764=>X"00",
1765=>X"00",
1766=>X"00",
1767=>X"00",
1768=>X"00",
1769=>X"00",
1770=>X"00",
1771=>X"00",
1772=>X"00",
1773=>X"00",
1774=>X"00",
1775=>X"00",
1776=>X"00",
1777=>X"00",
1778=>X"00",
1779=>X"00",
1780=>X"00",
1781=>X"00",
1782=>X"00",
1783=>X"00",
1784=>X"00",
1785=>X"00",
1786=>X"00",
1787=>X"00",
1788=>X"00",
1789=>X"00",
1790=>X"00",
1791=>X"00",
1792=>X"15",
1793=>X"15",
1794=>X"15",
1795=>X"15",
1796=>X"15",
1797=>X"15",
1798=>X"15",
1799=>X"15",
1800=>X"15",
1801=>X"15",
1802=>X"15",
1803=>X"15",
1804=>X"15",
1805=>X"15",
1806=>X"15",
1807=>X"15",
1808=>X"15",
1809=>X"15",
1810=>X"15",
1811=>X"15",
1812=>X"15",
1813=>X"15",
1814=>X"15",
1815=>X"15",
1816=>X"15",
1817=>X"15",
1818=>X"15",
1819=>X"15",
1820=>X"15",
1821=>X"15",
1822=>X"15",
1823=>X"15",
1824=>X"15",
1825=>X"15",
1826=>X"15",
1827=>X"15",
1828=>X"15",
1829=>X"15",
1830=>X"25",
1831=>X"15",
1832=>X"25",
1833=>X"15",
1834=>X"25",
1835=>X"15",
1836=>X"25",
1837=>X"25",
1838=>X"25",
1839=>X"25",
1840=>X"25",
1841=>X"25",
1842=>X"25",
1843=>X"25",
1844=>X"25",
1845=>X"25",
1846=>X"25",
1847=>X"25",
1848=>X"25",
1849=>X"25",
1850=>X"25",
1851=>X"25",
1852=>X"25",
1853=>X"25",
1854=>X"25",
1855=>X"25",
1856=>X"25",
1857=>X"15",
1858=>X"25",
1859=>X"15",
1860=>X"25",
1861=>X"25",
1862=>X"15",
1863=>X"25",
1864=>X"15",
1865=>X"25",
1866=>X"15",
1867=>X"25",
1868=>X"25",
1869=>X"15",
1870=>X"15",
1871=>X"25",
1872=>X"15",
1873=>X"15",
1874=>X"15",
1875=>X"15",
1876=>X"15",
1877=>X"15",
1878=>X"15",
1879=>X"15",
1880=>X"15",
1881=>X"15",
1882=>X"15",
1883=>X"15",
1884=>X"15",
1885=>X"15",
1886=>X"15",
1887=>X"15",
1888=>X"15",
1889=>X"15",
1890=>X"15",
1891=>X"15",
1892=>X"00",
1893=>X"00",
1894=>X"00",
1895=>X"00",
1896=>X"00",
1897=>X"00",
1898=>X"00",
1899=>X"00",
1900=>X"00",
1901=>X"00",
1902=>X"00",
1903=>X"00",
1904=>X"00",
1905=>X"00",
1906=>X"00",
1907=>X"00",
1908=>X"00",
1909=>X"00",
1910=>X"00",
1911=>X"00",
1912=>X"00",
1913=>X"00",
1914=>X"00",
1915=>X"00",
1916=>X"00",
1917=>X"00",
1918=>X"00",
1919=>X"00",
1920=>X"00",
1921=>X"00",
1922=>X"00",
1923=>X"00",
1924=>X"00",
1925=>X"00",
1926=>X"00",
1927=>X"00",
1928=>X"00",
1929=>X"00",
1930=>X"00",
1931=>X"00",
1932=>X"00",
1933=>X"00",
1934=>X"00",
1935=>X"00",
1936=>X"00",
1937=>X"00",
1938=>X"00",
1939=>X"00",
1940=>X"00",
1941=>X"00",
1942=>X"00",
1943=>X"00",
1944=>X"00",
1945=>X"00",
1946=>X"00",
1947=>X"00",
1948=>X"00",
1949=>X"00",
1950=>X"00",
1951=>X"00",
1952=>X"00",
1953=>X"00",
1954=>X"00",
1955=>X"00",
1956=>X"00",
1957=>X"00",
1958=>X"00",
1959=>X"00",
1960=>X"00",
1961=>X"00",
1962=>X"00",
1963=>X"00",
1964=>X"00",
1965=>X"00",
1966=>X"00",
1967=>X"00",
1968=>X"00",
1969=>X"00",
1970=>X"00",
1971=>X"00",
1972=>X"00",
1973=>X"00",
1974=>X"00",
1975=>X"00",
1976=>X"00",
1977=>X"00",
1978=>X"00",
1979=>X"00",
1980=>X"00",
1981=>X"00",
1982=>X"00",
1983=>X"00",
1984=>X"00",
1985=>X"00",
1986=>X"00",
1987=>X"00",
1988=>X"00",
1989=>X"00",
1990=>X"00",
1991=>X"00",
1992=>X"00",
1993=>X"00",
1994=>X"00",
1995=>X"00",
1996=>X"00",
1997=>X"00",
1998=>X"00",
1999=>X"00",
2000=>X"00",
2001=>X"00",
2002=>X"00",
2003=>X"00",
2004=>X"00",
2005=>X"00",
2006=>X"00",
2007=>X"00",
2008=>X"00",
2009=>X"00",
2010=>X"00",
2011=>X"00",
2012=>X"00",
2013=>X"00",
2014=>X"00",
2015=>X"00",
2016=>X"00",
2017=>X"00",
2018=>X"00",
2019=>X"00",
2020=>X"00",
2021=>X"00",
2022=>X"00",
2023=>X"00",
2024=>X"00",
2025=>X"00",
2026=>X"00",
2027=>X"00",
2028=>X"00",
2029=>X"00",
2030=>X"00",
2031=>X"00",
2032=>X"00",
2033=>X"00",
2034=>X"00",
2035=>X"00",
2036=>X"00",
2037=>X"00",
2038=>X"00",
2039=>X"00",
2040=>X"00",
2041=>X"00",
2042=>X"00",
2043=>X"00",
2044=>X"00",
2045=>X"00",
2046=>X"00",
2047=>X"00",
2048=>X"15",
2049=>X"15",
2050=>X"15",
2051=>X"15",
2052=>X"15",
2053=>X"15",
2054=>X"15",
2055=>X"15",
2056=>X"15",
2057=>X"15",
2058=>X"15",
2059=>X"15",
2060=>X"15",
2061=>X"15",
2062=>X"15",
2063=>X"15",
2064=>X"15",
2065=>X"15",
2066=>X"15",
2067=>X"15",
2068=>X"15",
2069=>X"15",
2070=>X"15",
2071=>X"15",
2072=>X"15",
2073=>X"15",
2074=>X"15",
2075=>X"15",
2076=>X"15",
2077=>X"15",
2078=>X"15",
2079=>X"15",
2080=>X"15",
2081=>X"15",
2082=>X"15",
2083=>X"15",
2084=>X"15",
2085=>X"25",
2086=>X"25",
2087=>X"15",
2088=>X"25",
2089=>X"15",
2090=>X"25",
2091=>X"15",
2092=>X"25",
2093=>X"25",
2094=>X"25",
2095=>X"25",
2096=>X"25",
2097=>X"25",
2098=>X"25",
2099=>X"25",
2100=>X"25",
2101=>X"25",
2102=>X"25",
2103=>X"25",
2104=>X"25",
2105=>X"25",
2106=>X"25",
2107=>X"25",
2108=>X"25",
2109=>X"25",
2110=>X"25",
2111=>X"25",
2112=>X"25",
2113=>X"15",
2114=>X"25",
2115=>X"15",
2116=>X"25",
2117=>X"25",
2118=>X"15",
2119=>X"25",
2120=>X"15",
2121=>X"25",
2122=>X"15",
2123=>X"25",
2124=>X"15",
2125=>X"25",
2126=>X"15",
2127=>X"25",
2128=>X"15",
2129=>X"15",
2130=>X"25",
2131=>X"15",
2132=>X"15",
2133=>X"15",
2134=>X"15",
2135=>X"15",
2136=>X"15",
2137=>X"15",
2138=>X"15",
2139=>X"15",
2140=>X"15",
2141=>X"15",
2142=>X"15",
2143=>X"15",
2144=>X"15",
2145=>X"15",
2146=>X"15",
2147=>X"15",
2148=>X"00",
2149=>X"00",
2150=>X"00",
2151=>X"00",
2152=>X"00",
2153=>X"00",
2154=>X"00",
2155=>X"00",
2156=>X"00",
2157=>X"00",
2158=>X"00",
2159=>X"00",
2160=>X"00",
2161=>X"00",
2162=>X"00",
2163=>X"00",
2164=>X"00",
2165=>X"00",
2166=>X"00",
2167=>X"00",
2168=>X"00",
2169=>X"00",
2170=>X"00",
2171=>X"00",
2172=>X"00",
2173=>X"00",
2174=>X"00",
2175=>X"00",
2176=>X"00",
2177=>X"00",
2178=>X"00",
2179=>X"00",
2180=>X"00",
2181=>X"00",
2182=>X"00",
2183=>X"00",
2184=>X"00",
2185=>X"00",
2186=>X"00",
2187=>X"00",
2188=>X"00",
2189=>X"00",
2190=>X"00",
2191=>X"00",
2192=>X"00",
2193=>X"00",
2194=>X"00",
2195=>X"00",
2196=>X"00",
2197=>X"00",
2198=>X"00",
2199=>X"00",
2200=>X"00",
2201=>X"00",
2202=>X"00",
2203=>X"00",
2204=>X"00",
2205=>X"00",
2206=>X"00",
2207=>X"00",
2208=>X"00",
2209=>X"00",
2210=>X"00",
2211=>X"00",
2212=>X"00",
2213=>X"00",
2214=>X"00",
2215=>X"00",
2216=>X"00",
2217=>X"00",
2218=>X"00",
2219=>X"00",
2220=>X"00",
2221=>X"00",
2222=>X"00",
2223=>X"00",
2224=>X"00",
2225=>X"00",
2226=>X"00",
2227=>X"00",
2228=>X"00",
2229=>X"00",
2230=>X"00",
2231=>X"00",
2232=>X"00",
2233=>X"00",
2234=>X"00",
2235=>X"00",
2236=>X"00",
2237=>X"00",
2238=>X"00",
2239=>X"00",
2240=>X"00",
2241=>X"00",
2242=>X"00",
2243=>X"00",
2244=>X"00",
2245=>X"00",
2246=>X"00",
2247=>X"00",
2248=>X"00",
2249=>X"00",
2250=>X"00",
2251=>X"00",
2252=>X"00",
2253=>X"00",
2254=>X"00",
2255=>X"00",
2256=>X"00",
2257=>X"00",
2258=>X"00",
2259=>X"00",
2260=>X"00",
2261=>X"00",
2262=>X"00",
2263=>X"00",
2264=>X"00",
2265=>X"00",
2266=>X"00",
2267=>X"00",
2268=>X"00",
2269=>X"00",
2270=>X"00",
2271=>X"00",
2272=>X"00",
2273=>X"00",
2274=>X"00",
2275=>X"00",
2276=>X"00",
2277=>X"00",
2278=>X"00",
2279=>X"00",
2280=>X"00",
2281=>X"00",
2282=>X"00",
2283=>X"00",
2284=>X"00",
2285=>X"00",
2286=>X"00",
2287=>X"00",
2288=>X"00",
2289=>X"00",
2290=>X"00",
2291=>X"00",
2292=>X"00",
2293=>X"00",
2294=>X"00",
2295=>X"00",
2296=>X"00",
2297=>X"00",
2298=>X"00",
2299=>X"00",
2300=>X"00",
2301=>X"00",
2302=>X"00",
2303=>X"00",
2304=>X"15",
2305=>X"15",
2306=>X"15",
2307=>X"15",
2308=>X"15",
2309=>X"15",
2310=>X"15",
2311=>X"15",
2312=>X"15",
2313=>X"15",
2314=>X"15",
2315=>X"15",
2316=>X"15",
2317=>X"15",
2318=>X"15",
2319=>X"15",
2320=>X"15",
2321=>X"15",
2322=>X"15",
2323=>X"15",
2324=>X"15",
2325=>X"15",
2326=>X"15",
2327=>X"15",
2328=>X"15",
2329=>X"15",
2330=>X"15",
2331=>X"15",
2332=>X"15",
2333=>X"15",
2334=>X"15",
2335=>X"15",
2336=>X"15",
2337=>X"15",
2338=>X"15",
2339=>X"15",
2340=>X"15",
2341=>X"25",
2342=>X"15",
2343=>X"15",
2344=>X"25",
2345=>X"15",
2346=>X"25",
2347=>X"15",
2348=>X"25",
2349=>X"15",
2350=>X"25",
2351=>X"15",
2352=>X"25",
2353=>X"25",
2354=>X"25",
2355=>X"25",
2356=>X"25",
2357=>X"25",
2358=>X"25",
2359=>X"25",
2360=>X"25",
2361=>X"25",
2362=>X"25",
2363=>X"25",
2364=>X"25",
2365=>X"25",
2366=>X"25",
2367=>X"25",
2368=>X"25",
2369=>X"25",
2370=>X"25",
2371=>X"25",
2372=>X"25",
2373=>X"25",
2374=>X"15",
2375=>X"25",
2376=>X"15",
2377=>X"25",
2378=>X"15",
2379=>X"25",
2380=>X"15",
2381=>X"25",
2382=>X"15",
2383=>X"15",
2384=>X"15",
2385=>X"15",
2386=>X"25",
2387=>X"15",
2388=>X"15",
2389=>X"15",
2390=>X"15",
2391=>X"15",
2392=>X"15",
2393=>X"15",
2394=>X"15",
2395=>X"15",
2396=>X"15",
2397=>X"19",
2398=>X"15",
2399=>X"15",
2400=>X"15",
2401=>X"15",
2402=>X"15",
2403=>X"15",
2404=>X"00",
2405=>X"00",
2406=>X"00",
2407=>X"00",
2408=>X"00",
2409=>X"00",
2410=>X"00",
2411=>X"00",
2412=>X"00",
2413=>X"00",
2414=>X"00",
2415=>X"00",
2416=>X"00",
2417=>X"00",
2418=>X"00",
2419=>X"00",
2420=>X"00",
2421=>X"00",
2422=>X"00",
2423=>X"00",
2424=>X"00",
2425=>X"00",
2426=>X"00",
2427=>X"00",
2428=>X"00",
2429=>X"00",
2430=>X"00",
2431=>X"00",
2432=>X"00",
2433=>X"00",
2434=>X"00",
2435=>X"00",
2436=>X"00",
2437=>X"00",
2438=>X"00",
2439=>X"00",
2440=>X"00",
2441=>X"00",
2442=>X"00",
2443=>X"00",
2444=>X"00",
2445=>X"00",
2446=>X"00",
2447=>X"00",
2448=>X"00",
2449=>X"00",
2450=>X"00",
2451=>X"00",
2452=>X"00",
2453=>X"00",
2454=>X"00",
2455=>X"00",
2456=>X"00",
2457=>X"00",
2458=>X"00",
2459=>X"00",
2460=>X"00",
2461=>X"00",
2462=>X"00",
2463=>X"00",
2464=>X"00",
2465=>X"00",
2466=>X"00",
2467=>X"00",
2468=>X"00",
2469=>X"00",
2470=>X"00",
2471=>X"00",
2472=>X"00",
2473=>X"00",
2474=>X"00",
2475=>X"00",
2476=>X"00",
2477=>X"00",
2478=>X"00",
2479=>X"00",
2480=>X"00",
2481=>X"00",
2482=>X"00",
2483=>X"00",
2484=>X"00",
2485=>X"00",
2486=>X"00",
2487=>X"00",
2488=>X"00",
2489=>X"00",
2490=>X"00",
2491=>X"00",
2492=>X"00",
2493=>X"00",
2494=>X"00",
2495=>X"00",
2496=>X"00",
2497=>X"00",
2498=>X"00",
2499=>X"00",
2500=>X"00",
2501=>X"00",
2502=>X"00",
2503=>X"00",
2504=>X"00",
2505=>X"00",
2506=>X"00",
2507=>X"00",
2508=>X"00",
2509=>X"00",
2510=>X"00",
2511=>X"00",
2512=>X"00",
2513=>X"00",
2514=>X"00",
2515=>X"00",
2516=>X"00",
2517=>X"00",
2518=>X"00",
2519=>X"00",
2520=>X"00",
2521=>X"00",
2522=>X"00",
2523=>X"00",
2524=>X"00",
2525=>X"00",
2526=>X"00",
2527=>X"00",
2528=>X"00",
2529=>X"00",
2530=>X"00",
2531=>X"00",
2532=>X"00",
2533=>X"00",
2534=>X"00",
2535=>X"00",
2536=>X"00",
2537=>X"00",
2538=>X"00",
2539=>X"00",
2540=>X"00",
2541=>X"00",
2542=>X"00",
2543=>X"00",
2544=>X"00",
2545=>X"00",
2546=>X"00",
2547=>X"00",
2548=>X"00",
2549=>X"00",
2550=>X"00",
2551=>X"00",
2552=>X"00",
2553=>X"00",
2554=>X"00",
2555=>X"00",
2556=>X"00",
2557=>X"00",
2558=>X"00",
2559=>X"00",
2560=>X"15",
2561=>X"15",
2562=>X"15",
2563=>X"15",
2564=>X"15",
2565=>X"15",
2566=>X"15",
2567=>X"15",
2568=>X"15",
2569=>X"15",
2570=>X"15",
2571=>X"15",
2572=>X"15",
2573=>X"15",
2574=>X"15",
2575=>X"15",
2576=>X"15",
2577=>X"15",
2578=>X"15",
2579=>X"15",
2580=>X"15",
2581=>X"15",
2582=>X"15",
2583=>X"15",
2584=>X"15",
2585=>X"15",
2586=>X"15",
2587=>X"15",
2588=>X"15",
2589=>X"15",
2590=>X"15",
2591=>X"15",
2592=>X"15",
2593=>X"15",
2594=>X"15",
2595=>X"15",
2596=>X"15",
2597=>X"15",
2598=>X"15",
2599=>X"15",
2600=>X"25",
2601=>X"15",
2602=>X"25",
2603=>X"15",
2604=>X"15",
2605=>X"15",
2606=>X"15",
2607=>X"25",
2608=>X"25",
2609=>X"25",
2610=>X"25",
2611=>X"25",
2612=>X"25",
2613=>X"25",
2614=>X"25",
2615=>X"25",
2616=>X"25",
2617=>X"25",
2618=>X"25",
2619=>X"25",
2620=>X"25",
2621=>X"25",
2622=>X"25",
2623=>X"25",
2624=>X"25",
2625=>X"25",
2626=>X"25",
2627=>X"25",
2628=>X"15",
2629=>X"15",
2630=>X"15",
2631=>X"15",
2632=>X"25",
2633=>X"25",
2634=>X"15",
2635=>X"25",
2636=>X"15",
2637=>X"15",
2638=>X"15",
2639=>X"15",
2640=>X"15",
2641=>X"15",
2642=>X"15",
2643=>X"15",
2644=>X"15",
2645=>X"15",
2646=>X"15",
2647=>X"15",
2648=>X"15",
2649=>X"15",
2650=>X"15",
2651=>X"15",
2652=>X"15",
2653=>X"19",
2654=>X"15",
2655=>X"15",
2656=>X"15",
2657=>X"15",
2658=>X"15",
2659=>X"15",
2660=>X"00",
2661=>X"00",
2662=>X"00",
2663=>X"00",
2664=>X"00",
2665=>X"00",
2666=>X"00",
2667=>X"00",
2668=>X"00",
2669=>X"00",
2670=>X"00",
2671=>X"00",
2672=>X"00",
2673=>X"00",
2674=>X"00",
2675=>X"00",
2676=>X"00",
2677=>X"00",
2678=>X"00",
2679=>X"00",
2680=>X"00",
2681=>X"00",
2682=>X"00",
2683=>X"00",
2684=>X"00",
2685=>X"00",
2686=>X"00",
2687=>X"00",
2688=>X"00",
2689=>X"00",
2690=>X"00",
2691=>X"00",
2692=>X"00",
2693=>X"00",
2694=>X"00",
2695=>X"00",
2696=>X"00",
2697=>X"00",
2698=>X"00",
2699=>X"00",
2700=>X"00",
2701=>X"00",
2702=>X"00",
2703=>X"00",
2704=>X"00",
2705=>X"00",
2706=>X"00",
2707=>X"00",
2708=>X"00",
2709=>X"00",
2710=>X"00",
2711=>X"00",
2712=>X"00",
2713=>X"00",
2714=>X"00",
2715=>X"00",
2716=>X"00",
2717=>X"00",
2718=>X"00",
2719=>X"00",
2720=>X"00",
2721=>X"00",
2722=>X"00",
2723=>X"00",
2724=>X"00",
2725=>X"00",
2726=>X"00",
2727=>X"00",
2728=>X"00",
2729=>X"00",
2730=>X"00",
2731=>X"00",
2732=>X"00",
2733=>X"00",
2734=>X"00",
2735=>X"00",
2736=>X"00",
2737=>X"00",
2738=>X"00",
2739=>X"00",
2740=>X"00",
2741=>X"00",
2742=>X"00",
2743=>X"00",
2744=>X"00",
2745=>X"00",
2746=>X"00",
2747=>X"00",
2748=>X"00",
2749=>X"00",
2750=>X"00",
2751=>X"00",
2752=>X"00",
2753=>X"00",
2754=>X"00",
2755=>X"00",
2756=>X"00",
2757=>X"00",
2758=>X"00",
2759=>X"00",
2760=>X"00",
2761=>X"00",
2762=>X"00",
2763=>X"00",
2764=>X"00",
2765=>X"00",
2766=>X"00",
2767=>X"00",
2768=>X"00",
2769=>X"00",
2770=>X"00",
2771=>X"00",
2772=>X"00",
2773=>X"00",
2774=>X"00",
2775=>X"00",
2776=>X"00",
2777=>X"00",
2778=>X"00",
2779=>X"00",
2780=>X"00",
2781=>X"00",
2782=>X"00",
2783=>X"00",
2784=>X"00",
2785=>X"00",
2786=>X"00",
2787=>X"00",
2788=>X"00",
2789=>X"00",
2790=>X"00",
2791=>X"00",
2792=>X"00",
2793=>X"00",
2794=>X"00",
2795=>X"00",
2796=>X"00",
2797=>X"00",
2798=>X"00",
2799=>X"00",
2800=>X"00",
2801=>X"00",
2802=>X"00",
2803=>X"00",
2804=>X"00",
2805=>X"00",
2806=>X"00",
2807=>X"00",
2808=>X"00",
2809=>X"00",
2810=>X"00",
2811=>X"00",
2812=>X"00",
2813=>X"00",
2814=>X"00",
2815=>X"00",
2816=>X"15",
2817=>X"15",
2818=>X"15",
2819=>X"15",
2820=>X"15",
2821=>X"15",
2822=>X"15",
2823=>X"15",
2824=>X"15",
2825=>X"15",
2826=>X"15",
2827=>X"15",
2828=>X"15",
2829=>X"15",
2830=>X"15",
2831=>X"15",
2832=>X"15",
2833=>X"15",
2834=>X"15",
2835=>X"15",
2836=>X"15",
2837=>X"15",
2838=>X"15",
2839=>X"15",
2840=>X"15",
2841=>X"15",
2842=>X"15",
2843=>X"25",
2844=>X"15",
2845=>X"15",
2846=>X"25",
2847=>X"15",
2848=>X"25",
2849=>X"15",
2850=>X"15",
2851=>X"25",
2852=>X"15",
2853=>X"25",
2854=>X"15",
2855=>X"25",
2856=>X"15",
2857=>X"15",
2858=>X"15",
2859=>X"15",
2860=>X"15",
2861=>X"25",
2862=>X"25",
2863=>X"25",
2864=>X"25",
2865=>X"25",
2866=>X"25",
2867=>X"25",
2868=>X"25",
2869=>X"29",
2870=>X"25",
2871=>X"25",
2872=>X"25",
2873=>X"25",
2874=>X"25",
2875=>X"25",
2876=>X"25",
2877=>X"25",
2878=>X"25",
2879=>X"25",
2880=>X"25",
2881=>X"25",
2882=>X"25",
2883=>X"25",
2884=>X"25",
2885=>X"25",
2886=>X"15",
2887=>X"25",
2888=>X"25",
2889=>X"25",
2890=>X"15",
2891=>X"25",
2892=>X"15",
2893=>X"25",
2894=>X"15",
2895=>X"25",
2896=>X"15",
2897=>X"15",
2898=>X"15",
2899=>X"15",
2900=>X"25",
2901=>X"15",
2902=>X"15",
2903=>X"15",
2904=>X"15",
2905=>X"15",
2906=>X"15",
2907=>X"29",
2908=>X"15",
2909=>X"15",
2910=>X"15",
2911=>X"15",
2912=>X"15",
2913=>X"15",
2914=>X"15",
2915=>X"15",
2916=>X"00",
2917=>X"00",
2918=>X"00",
2919=>X"00",
2920=>X"00",
2921=>X"00",
2922=>X"00",
2923=>X"00",
2924=>X"00",
2925=>X"00",
2926=>X"00",
2927=>X"00",
2928=>X"00",
2929=>X"00",
2930=>X"00",
2931=>X"00",
2932=>X"00",
2933=>X"00",
2934=>X"00",
2935=>X"00",
2936=>X"00",
2937=>X"00",
2938=>X"00",
2939=>X"00",
2940=>X"00",
2941=>X"00",
2942=>X"00",
2943=>X"00",
2944=>X"00",
2945=>X"00",
2946=>X"00",
2947=>X"00",
2948=>X"00",
2949=>X"00",
2950=>X"00",
2951=>X"00",
2952=>X"00",
2953=>X"00",
2954=>X"00",
2955=>X"00",
2956=>X"00",
2957=>X"00",
2958=>X"00",
2959=>X"00",
2960=>X"00",
2961=>X"00",
2962=>X"00",
2963=>X"00",
2964=>X"00",
2965=>X"00",
2966=>X"00",
2967=>X"00",
2968=>X"00",
2969=>X"00",
2970=>X"00",
2971=>X"00",
2972=>X"00",
2973=>X"00",
2974=>X"00",
2975=>X"00",
2976=>X"00",
2977=>X"00",
2978=>X"00",
2979=>X"00",
2980=>X"00",
2981=>X"00",
2982=>X"00",
2983=>X"00",
2984=>X"00",
2985=>X"00",
2986=>X"00",
2987=>X"00",
2988=>X"00",
2989=>X"00",
2990=>X"00",
2991=>X"00",
2992=>X"00",
2993=>X"00",
2994=>X"00",
2995=>X"00",
2996=>X"00",
2997=>X"00",
2998=>X"00",
2999=>X"00",
3000=>X"00",
3001=>X"00",
3002=>X"00",
3003=>X"00",
3004=>X"00",
3005=>X"00",
3006=>X"00",
3007=>X"00",
3008=>X"00",
3009=>X"00",
3010=>X"00",
3011=>X"00",
3012=>X"00",
3013=>X"00",
3014=>X"00",
3015=>X"00",
3016=>X"00",
3017=>X"00",
3018=>X"00",
3019=>X"00",
3020=>X"00",
3021=>X"00",
3022=>X"00",
3023=>X"00",
3024=>X"00",
3025=>X"00",
3026=>X"00",
3027=>X"00",
3028=>X"00",
3029=>X"00",
3030=>X"00",
3031=>X"00",
3032=>X"00",
3033=>X"00",
3034=>X"00",
3035=>X"00",
3036=>X"00",
3037=>X"00",
3038=>X"00",
3039=>X"00",
3040=>X"00",
3041=>X"00",
3042=>X"00",
3043=>X"00",
3044=>X"00",
3045=>X"00",
3046=>X"00",
3047=>X"00",
3048=>X"00",
3049=>X"00",
3050=>X"00",
3051=>X"00",
3052=>X"00",
3053=>X"00",
3054=>X"00",
3055=>X"00",
3056=>X"00",
3057=>X"00",
3058=>X"00",
3059=>X"00",
3060=>X"00",
3061=>X"00",
3062=>X"00",
3063=>X"00",
3064=>X"00",
3065=>X"00",
3066=>X"00",
3067=>X"00",
3068=>X"00",
3069=>X"00",
3070=>X"00",
3071=>X"00",
3072=>X"15",
3073=>X"15",
3074=>X"15",
3075=>X"15",
3076=>X"15",
3077=>X"15",
3078=>X"15",
3079=>X"15",
3080=>X"15",
3081=>X"15",
3082=>X"15",
3083=>X"15",
3084=>X"15",
3085=>X"15",
3086=>X"15",
3087=>X"15",
3088=>X"15",
3089=>X"15",
3090=>X"15",
3091=>X"15",
3092=>X"15",
3093=>X"15",
3094=>X"15",
3095=>X"15",
3096=>X"15",
3097=>X"15",
3098=>X"25",
3099=>X"25",
3100=>X"15",
3101=>X"15",
3102=>X"25",
3103=>X"25",
3104=>X"15",
3105=>X"15",
3106=>X"25",
3107=>X"25",
3108=>X"15",
3109=>X"15",
3110=>X"25",
3111=>X"25",
3112=>X"15",
3113=>X"15",
3114=>X"15",
3115=>X"15",
3116=>X"15",
3117=>X"15",
3118=>X"25",
3119=>X"25",
3120=>X"15",
3121=>X"15",
3122=>X"25",
3123=>X"25",
3124=>X"29",
3125=>X"29",
3126=>X"25",
3127=>X"25",
3128=>X"25",
3129=>X"25",
3130=>X"25",
3131=>X"25",
3132=>X"25",
3133=>X"25",
3134=>X"25",
3135=>X"25",
3136=>X"25",
3137=>X"25",
3138=>X"25",
3139=>X"25",
3140=>X"25",
3141=>X"25",
3142=>X"25",
3143=>X"15",
3144=>X"25",
3145=>X"25",
3146=>X"25",
3147=>X"25",
3148=>X"25",
3149=>X"25",
3150=>X"15",
3151=>X"15",
3152=>X"15",
3153=>X"15",
3154=>X"15",
3155=>X"15",
3156=>X"15",
3157=>X"15",
3158=>X"15",
3159=>X"15",
3160=>X"15",
3161=>X"15",
3162=>X"25",
3163=>X"25",
3164=>X"15",
3165=>X"15",
3166=>X"15",
3167=>X"15",
3168=>X"15",
3169=>X"15",
3170=>X"15",
3171=>X"15",
3172=>X"00",
3173=>X"00",
3174=>X"00",
3175=>X"00",
3176=>X"00",
3177=>X"00",
3178=>X"00",
3179=>X"00",
3180=>X"00",
3181=>X"00",
3182=>X"00",
3183=>X"00",
3184=>X"00",
3185=>X"00",
3186=>X"00",
3187=>X"00",
3188=>X"00",
3189=>X"00",
3190=>X"00",
3191=>X"00",
3192=>X"00",
3193=>X"00",
3194=>X"00",
3195=>X"00",
3196=>X"00",
3197=>X"00",
3198=>X"00",
3199=>X"00",
3200=>X"00",
3201=>X"00",
3202=>X"00",
3203=>X"00",
3204=>X"00",
3205=>X"00",
3206=>X"00",
3207=>X"00",
3208=>X"00",
3209=>X"00",
3210=>X"00",
3211=>X"00",
3212=>X"00",
3213=>X"00",
3214=>X"00",
3215=>X"00",
3216=>X"00",
3217=>X"00",
3218=>X"00",
3219=>X"00",
3220=>X"00",
3221=>X"00",
3222=>X"00",
3223=>X"00",
3224=>X"00",
3225=>X"00",
3226=>X"00",
3227=>X"00",
3228=>X"00",
3229=>X"00",
3230=>X"00",
3231=>X"00",
3232=>X"00",
3233=>X"00",
3234=>X"00",
3235=>X"00",
3236=>X"00",
3237=>X"00",
3238=>X"00",
3239=>X"00",
3240=>X"00",
3241=>X"00",
3242=>X"00",
3243=>X"00",
3244=>X"00",
3245=>X"00",
3246=>X"00",
3247=>X"00",
3248=>X"00",
3249=>X"00",
3250=>X"00",
3251=>X"00",
3252=>X"00",
3253=>X"00",
3254=>X"00",
3255=>X"00",
3256=>X"00",
3257=>X"00",
3258=>X"00",
3259=>X"00",
3260=>X"00",
3261=>X"00",
3262=>X"00",
3263=>X"00",
3264=>X"00",
3265=>X"00",
3266=>X"00",
3267=>X"00",
3268=>X"00",
3269=>X"00",
3270=>X"00",
3271=>X"00",
3272=>X"00",
3273=>X"00",
3274=>X"00",
3275=>X"00",
3276=>X"00",
3277=>X"00",
3278=>X"00",
3279=>X"00",
3280=>X"00",
3281=>X"00",
3282=>X"00",
3283=>X"00",
3284=>X"00",
3285=>X"00",
3286=>X"00",
3287=>X"00",
3288=>X"00",
3289=>X"00",
3290=>X"00",
3291=>X"00",
3292=>X"00",
3293=>X"00",
3294=>X"00",
3295=>X"00",
3296=>X"00",
3297=>X"00",
3298=>X"00",
3299=>X"00",
3300=>X"00",
3301=>X"00",
3302=>X"00",
3303=>X"00",
3304=>X"00",
3305=>X"00",
3306=>X"00",
3307=>X"00",
3308=>X"00",
3309=>X"00",
3310=>X"00",
3311=>X"00",
3312=>X"00",
3313=>X"00",
3314=>X"00",
3315=>X"00",
3316=>X"00",
3317=>X"00",
3318=>X"00",
3319=>X"00",
3320=>X"00",
3321=>X"00",
3322=>X"00",
3323=>X"00",
3324=>X"00",
3325=>X"00",
3326=>X"00",
3327=>X"00",
3328=>X"15",
3329=>X"15",
3330=>X"15",
3331=>X"15",
3332=>X"15",
3333=>X"15",
3334=>X"15",
3335=>X"15",
3336=>X"15",
3337=>X"15",
3338=>X"15",
3339=>X"15",
3340=>X"15",
3341=>X"15",
3342=>X"15",
3343=>X"15",
3344=>X"15",
3345=>X"15",
3346=>X"15",
3347=>X"15",
3348=>X"15",
3349=>X"15",
3350=>X"15",
3351=>X"15",
3352=>X"15",
3353=>X"15",
3354=>X"15",
3355=>X"15",
3356=>X"15",
3357=>X"15",
3358=>X"15",
3359=>X"15",
3360=>X"15",
3361=>X"15",
3362=>X"15",
3363=>X"15",
3364=>X"15",
3365=>X"25",
3366=>X"15",
3367=>X"15",
3368=>X"15",
3369=>X"25",
3370=>X"15",
3371=>X"15",
3372=>X"25",
3373=>X"15",
3374=>X"15",
3375=>X"15",
3376=>X"25",
3377=>X"25",
3378=>X"15",
3379=>X"29",
3380=>X"25",
3381=>X"25",
3382=>X"2A",
3383=>X"2A",
3384=>X"29",
3385=>X"29",
3386=>X"35",
3387=>X"35",
3388=>X"25",
3389=>X"25",
3390=>X"25",
3391=>X"25",
3392=>X"25",
3393=>X"25",
3394=>X"25",
3395=>X"25",
3396=>X"25",
3397=>X"25",
3398=>X"25",
3399=>X"25",
3400=>X"15",
3401=>X"25",
3402=>X"25",
3403=>X"15",
3404=>X"15",
3405=>X"15",
3406=>X"15",
3407=>X"15",
3408=>X"25",
3409=>X"15",
3410=>X"15",
3411=>X"15",
3412=>X"15",
3413=>X"19",
3414=>X"15",
3415=>X"25",
3416=>X"15",
3417=>X"15",
3418=>X"15",
3419=>X"15",
3420=>X"15",
3421=>X"15",
3422=>X"15",
3423=>X"15",
3424=>X"15",
3425=>X"15",
3426=>X"15",
3427=>X"15",
3428=>X"00",
3429=>X"00",
3430=>X"00",
3431=>X"00",
3432=>X"00",
3433=>X"00",
3434=>X"00",
3435=>X"00",
3436=>X"00",
3437=>X"00",
3438=>X"00",
3439=>X"00",
3440=>X"00",
3441=>X"00",
3442=>X"00",
3443=>X"00",
3444=>X"00",
3445=>X"00",
3446=>X"00",
3447=>X"00",
3448=>X"00",
3449=>X"00",
3450=>X"00",
3451=>X"00",
3452=>X"00",
3453=>X"00",
3454=>X"00",
3455=>X"00",
3456=>X"00",
3457=>X"00",
3458=>X"00",
3459=>X"00",
3460=>X"00",
3461=>X"00",
3462=>X"00",
3463=>X"00",
3464=>X"00",
3465=>X"00",
3466=>X"00",
3467=>X"00",
3468=>X"00",
3469=>X"00",
3470=>X"00",
3471=>X"00",
3472=>X"00",
3473=>X"00",
3474=>X"00",
3475=>X"00",
3476=>X"00",
3477=>X"00",
3478=>X"00",
3479=>X"00",
3480=>X"00",
3481=>X"00",
3482=>X"00",
3483=>X"00",
3484=>X"00",
3485=>X"00",
3486=>X"00",
3487=>X"00",
3488=>X"00",
3489=>X"00",
3490=>X"00",
3491=>X"00",
3492=>X"00",
3493=>X"00",
3494=>X"00",
3495=>X"00",
3496=>X"00",
3497=>X"00",
3498=>X"00",
3499=>X"00",
3500=>X"00",
3501=>X"00",
3502=>X"00",
3503=>X"00",
3504=>X"00",
3505=>X"00",
3506=>X"00",
3507=>X"00",
3508=>X"00",
3509=>X"00",
3510=>X"00",
3511=>X"00",
3512=>X"00",
3513=>X"00",
3514=>X"00",
3515=>X"00",
3516=>X"00",
3517=>X"00",
3518=>X"00",
3519=>X"00",
3520=>X"00",
3521=>X"00",
3522=>X"00",
3523=>X"00",
3524=>X"00",
3525=>X"00",
3526=>X"00",
3527=>X"00",
3528=>X"00",
3529=>X"00",
3530=>X"00",
3531=>X"00",
3532=>X"00",
3533=>X"00",
3534=>X"00",
3535=>X"00",
3536=>X"00",
3537=>X"00",
3538=>X"00",
3539=>X"00",
3540=>X"00",
3541=>X"00",
3542=>X"00",
3543=>X"00",
3544=>X"00",
3545=>X"00",
3546=>X"00",
3547=>X"00",
3548=>X"00",
3549=>X"00",
3550=>X"00",
3551=>X"00",
3552=>X"00",
3553=>X"00",
3554=>X"00",
3555=>X"00",
3556=>X"00",
3557=>X"00",
3558=>X"00",
3559=>X"00",
3560=>X"00",
3561=>X"00",
3562=>X"00",
3563=>X"00",
3564=>X"00",
3565=>X"00",
3566=>X"00",
3567=>X"00",
3568=>X"00",
3569=>X"00",
3570=>X"00",
3571=>X"00",
3572=>X"00",
3573=>X"00",
3574=>X"00",
3575=>X"00",
3576=>X"00",
3577=>X"00",
3578=>X"00",
3579=>X"00",
3580=>X"00",
3581=>X"00",
3582=>X"00",
3583=>X"00",
3584=>X"15",
3585=>X"15",
3586=>X"15",
3587=>X"15",
3588=>X"15",
3589=>X"15",
3590=>X"15",
3591=>X"15",
3592=>X"15",
3593=>X"15",
3594=>X"15",
3595=>X"15",
3596=>X"15",
3597=>X"15",
3598=>X"15",
3599=>X"15",
3600=>X"15",
3601=>X"15",
3602=>X"15",
3603=>X"15",
3604=>X"15",
3605=>X"15",
3606=>X"15",
3607=>X"15",
3608=>X"15",
3609=>X"15",
3610=>X"15",
3611=>X"15",
3612=>X"15",
3613=>X"15",
3614=>X"15",
3615=>X"15",
3616=>X"15",
3617=>X"15",
3618=>X"15",
3619=>X"15",
3620=>X"15",
3621=>X"15",
3622=>X"15",
3623=>X"15",
3624=>X"15",
3625=>X"15",
3626=>X"15",
3627=>X"15",
3628=>X"15",
3629=>X"15",
3630=>X"25",
3631=>X"15",
3632=>X"29",
3633=>X"25",
3634=>X"15",
3635=>X"15",
3636=>X"15",
3637=>X"2A",
3638=>X"2A",
3639=>X"2A",
3640=>X"2A",
3641=>X"39",
3642=>X"35",
3643=>X"39",
3644=>X"35",
3645=>X"25",
3646=>X"25",
3647=>X"25",
3648=>X"25",
3649=>X"25",
3650=>X"25",
3651=>X"25",
3652=>X"25",
3653=>X"25",
3654=>X"15",
3655=>X"25",
3656=>X"25",
3657=>X"15",
3658=>X"15",
3659=>X"25",
3660=>X"25",
3661=>X"15",
3662=>X"25",
3663=>X"15",
3664=>X"15",
3665=>X"15",
3666=>X"15",
3667=>X"15",
3668=>X"15",
3669=>X"15",
3670=>X"15",
3671=>X"15",
3672=>X"15",
3673=>X"15",
3674=>X"15",
3675=>X"15",
3676=>X"19",
3677=>X"15",
3678=>X"15",
3679=>X"15",
3680=>X"15",
3681=>X"15",
3682=>X"15",
3683=>X"15",
3684=>X"00",
3685=>X"00",
3686=>X"00",
3687=>X"00",
3688=>X"00",
3689=>X"00",
3690=>X"00",
3691=>X"00",
3692=>X"00",
3693=>X"00",
3694=>X"00",
3695=>X"00",
3696=>X"00",
3697=>X"00",
3698=>X"00",
3699=>X"00",
3700=>X"00",
3701=>X"00",
3702=>X"00",
3703=>X"00",
3704=>X"00",
3705=>X"00",
3706=>X"00",
3707=>X"00",
3708=>X"00",
3709=>X"00",
3710=>X"00",
3711=>X"00",
3712=>X"00",
3713=>X"00",
3714=>X"00",
3715=>X"00",
3716=>X"00",
3717=>X"00",
3718=>X"00",
3719=>X"00",
3720=>X"00",
3721=>X"00",
3722=>X"00",
3723=>X"00",
3724=>X"00",
3725=>X"00",
3726=>X"00",
3727=>X"00",
3728=>X"00",
3729=>X"00",
3730=>X"00",
3731=>X"00",
3732=>X"00",
3733=>X"00",
3734=>X"00",
3735=>X"00",
3736=>X"00",
3737=>X"00",
3738=>X"00",
3739=>X"00",
3740=>X"00",
3741=>X"00",
3742=>X"00",
3743=>X"00",
3744=>X"00",
3745=>X"00",
3746=>X"00",
3747=>X"00",
3748=>X"00",
3749=>X"00",
3750=>X"00",
3751=>X"00",
3752=>X"00",
3753=>X"00",
3754=>X"00",
3755=>X"00",
3756=>X"00",
3757=>X"00",
3758=>X"00",
3759=>X"00",
3760=>X"00",
3761=>X"00",
3762=>X"00",
3763=>X"00",
3764=>X"00",
3765=>X"00",
3766=>X"00",
3767=>X"00",
3768=>X"00",
3769=>X"00",
3770=>X"00",
3771=>X"00",
3772=>X"00",
3773=>X"00",
3774=>X"00",
3775=>X"00",
3776=>X"00",
3777=>X"00",
3778=>X"00",
3779=>X"00",
3780=>X"00",
3781=>X"00",
3782=>X"00",
3783=>X"00",
3784=>X"00",
3785=>X"00",
3786=>X"00",
3787=>X"00",
3788=>X"00",
3789=>X"00",
3790=>X"00",
3791=>X"00",
3792=>X"00",
3793=>X"00",
3794=>X"00",
3795=>X"00",
3796=>X"00",
3797=>X"00",
3798=>X"00",
3799=>X"00",
3800=>X"00",
3801=>X"00",
3802=>X"00",
3803=>X"00",
3804=>X"00",
3805=>X"00",
3806=>X"00",
3807=>X"00",
3808=>X"00",
3809=>X"00",
3810=>X"00",
3811=>X"00",
3812=>X"00",
3813=>X"00",
3814=>X"00",
3815=>X"00",
3816=>X"00",
3817=>X"00",
3818=>X"00",
3819=>X"00",
3820=>X"00",
3821=>X"00",
3822=>X"00",
3823=>X"00",
3824=>X"00",
3825=>X"00",
3826=>X"00",
3827=>X"00",
3828=>X"00",
3829=>X"00",
3830=>X"00",
3831=>X"00",
3832=>X"00",
3833=>X"00",
3834=>X"00",
3835=>X"00",
3836=>X"00",
3837=>X"00",
3838=>X"00",
3839=>X"00",
3840=>X"15",
3841=>X"15",
3842=>X"15",
3843=>X"15",
3844=>X"15",
3845=>X"15",
3846=>X"15",
3847=>X"15",
3848=>X"15",
3849=>X"15",
3850=>X"15",
3851=>X"15",
3852=>X"15",
3853=>X"15",
3854=>X"15",
3855=>X"15",
3856=>X"15",
3857=>X"15",
3858=>X"15",
3859=>X"15",
3860=>X"15",
3861=>X"15",
3862=>X"15",
3863=>X"15",
3864=>X"15",
3865=>X"15",
3866=>X"15",
3867=>X"15",
3868=>X"15",
3869=>X"15",
3870=>X"15",
3871=>X"15",
3872=>X"25",
3873=>X"15",
3874=>X"15",
3875=>X"15",
3876=>X"15",
3877=>X"15",
3878=>X"15",
3879=>X"25",
3880=>X"15",
3881=>X"15",
3882=>X"19",
3883=>X"15",
3884=>X"15",
3885=>X"15",
3886=>X"19",
3887=>X"15",
3888=>X"15",
3889=>X"15",
3890=>X"15",
3891=>X"19",
3892=>X"2E",
3893=>X"2F",
3894=>X"2F",
3895=>X"1F",
3896=>X"1F",
3897=>X"2B",
3898=>X"36",
3899=>X"35",
3900=>X"34",
3901=>X"35",
3902=>X"25",
3903=>X"25",
3904=>X"25",
3905=>X"25",
3906=>X"25",
3907=>X"25",
3908=>X"25",
3909=>X"25",
3910=>X"25",
3911=>X"25",
3912=>X"25",
3913=>X"25",
3914=>X"15",
3915=>X"25",
3916=>X"25",
3917=>X"15",
3918=>X"15",
3919=>X"15",
3920=>X"25",
3921=>X"15",
3922=>X"15",
3923=>X"25",
3924=>X"15",
3925=>X"15",
3926=>X"15",
3927=>X"15",
3928=>X"19",
3929=>X"15",
3930=>X"15",
3931=>X"15",
3932=>X"15",
3933=>X"15",
3934=>X"15",
3935=>X"15",
3936=>X"15",
3937=>X"15",
3938=>X"15",
3939=>X"15",
3940=>X"00",
3941=>X"00",
3942=>X"00",
3943=>X"00",
3944=>X"00",
3945=>X"00",
3946=>X"00",
3947=>X"00",
3948=>X"00",
3949=>X"00",
3950=>X"00",
3951=>X"00",
3952=>X"00",
3953=>X"00",
3954=>X"00",
3955=>X"00",
3956=>X"00",
3957=>X"00",
3958=>X"00",
3959=>X"00",
3960=>X"00",
3961=>X"00",
3962=>X"00",
3963=>X"00",
3964=>X"00",
3965=>X"00",
3966=>X"00",
3967=>X"00",
3968=>X"00",
3969=>X"00",
3970=>X"00",
3971=>X"00",
3972=>X"00",
3973=>X"00",
3974=>X"00",
3975=>X"00",
3976=>X"00",
3977=>X"00",
3978=>X"00",
3979=>X"00",
3980=>X"00",
3981=>X"00",
3982=>X"00",
3983=>X"00",
3984=>X"00",
3985=>X"00",
3986=>X"00",
3987=>X"00",
3988=>X"00",
3989=>X"00",
3990=>X"00",
3991=>X"00",
3992=>X"00",
3993=>X"00",
3994=>X"00",
3995=>X"00",
3996=>X"00",
3997=>X"00",
3998=>X"00",
3999=>X"00",
4000=>X"00",
4001=>X"00",
4002=>X"00",
4003=>X"00",
4004=>X"00",
4005=>X"00",
4006=>X"00",
4007=>X"00",
4008=>X"00",
4009=>X"00",
4010=>X"00",
4011=>X"00",
4012=>X"00",
4013=>X"00",
4014=>X"00",
4015=>X"00",
4016=>X"00",
4017=>X"00",
4018=>X"00",
4019=>X"00",
4020=>X"00",
4021=>X"00",
4022=>X"00",
4023=>X"00",
4024=>X"00",
4025=>X"00",
4026=>X"00",
4027=>X"00",
4028=>X"00",
4029=>X"00",
4030=>X"00",
4031=>X"00",
4032=>X"00",
4033=>X"00",
4034=>X"00",
4035=>X"00",
4036=>X"00",
4037=>X"00",
4038=>X"00",
4039=>X"00",
4040=>X"00",
4041=>X"00",
4042=>X"00",
4043=>X"00",
4044=>X"00",
4045=>X"00",
4046=>X"00",
4047=>X"00",
4048=>X"00",
4049=>X"00",
4050=>X"00",
4051=>X"00",
4052=>X"00",
4053=>X"00",
4054=>X"00",
4055=>X"00",
4056=>X"00",
4057=>X"00",
4058=>X"00",
4059=>X"00",
4060=>X"00",
4061=>X"00",
4062=>X"00",
4063=>X"00",
4064=>X"00",
4065=>X"00",
4066=>X"00",
4067=>X"00",
4068=>X"00",
4069=>X"00",
4070=>X"00",
4071=>X"00",
4072=>X"00",
4073=>X"00",
4074=>X"00",
4075=>X"00",
4076=>X"00",
4077=>X"00",
4078=>X"00",
4079=>X"00",
4080=>X"00",
4081=>X"00",
4082=>X"00",
4083=>X"00",
4084=>X"00",
4085=>X"00",
4086=>X"00",
4087=>X"00",
4088=>X"00",
4089=>X"00",
4090=>X"00",
4091=>X"00",
4092=>X"00",
4093=>X"00",
4094=>X"00",
4095=>X"00",
4096=>X"15",
4097=>X"15",
4098=>X"15",
4099=>X"15",
4100=>X"15",
4101=>X"15",
4102=>X"15",
4103=>X"15",
4104=>X"15",
4105=>X"15",
4106=>X"15",
4107=>X"15",
4108=>X"15",
4109=>X"15",
4110=>X"15",
4111=>X"15",
4112=>X"15",
4113=>X"15",
4114=>X"15",
4115=>X"15",
4116=>X"15",
4117=>X"15",
4118=>X"15",
4119=>X"15",
4120=>X"15",
4121=>X"15",
4122=>X"15",
4123=>X"15",
4124=>X"15",
4125=>X"15",
4126=>X"15",
4127=>X"15",
4128=>X"15",
4129=>X"15",
4130=>X"15",
4131=>X"15",
4132=>X"15",
4133=>X"19",
4134=>X"15",
4135=>X"19",
4136=>X"15",
4137=>X"15",
4138=>X"15",
4139=>X"15",
4140=>X"19",
4141=>X"15",
4142=>X"15",
4143=>X"15",
4144=>X"15",
4145=>X"29",
4146=>X"29",
4147=>X"2D",
4148=>X"3D",
4149=>X"2E",
4150=>X"2F",
4151=>X"1F",
4152=>X"1B",
4153=>X"1B",
4154=>X"2B",
4155=>X"35",
4156=>X"34",
4157=>X"34",
4158=>X"35",
4159=>X"35",
4160=>X"25",
4161=>X"25",
4162=>X"25",
4163=>X"25",
4164=>X"25",
4165=>X"25",
4166=>X"25",
4167=>X"25",
4168=>X"25",
4169=>X"25",
4170=>X"15",
4171=>X"15",
4172=>X"15",
4173=>X"15",
4174=>X"15",
4175=>X"15",
4176=>X"15",
4177=>X"15",
4178=>X"15",
4179=>X"15",
4180=>X"15",
4181=>X"15",
4182=>X"15",
4183=>X"15",
4184=>X"15",
4185=>X"15",
4186=>X"15",
4187=>X"15",
4188=>X"15",
4189=>X"15",
4190=>X"15",
4191=>X"15",
4192=>X"15",
4193=>X"15",
4194=>X"15",
4195=>X"15",
4196=>X"00",
4197=>X"00",
4198=>X"00",
4199=>X"00",
4200=>X"00",
4201=>X"00",
4202=>X"00",
4203=>X"00",
4204=>X"00",
4205=>X"00",
4206=>X"00",
4207=>X"00",
4208=>X"00",
4209=>X"00",
4210=>X"00",
4211=>X"00",
4212=>X"00",
4213=>X"00",
4214=>X"00",
4215=>X"00",
4216=>X"00",
4217=>X"00",
4218=>X"00",
4219=>X"00",
4220=>X"00",
4221=>X"00",
4222=>X"00",
4223=>X"00",
4224=>X"00",
4225=>X"00",
4226=>X"00",
4227=>X"00",
4228=>X"00",
4229=>X"00",
4230=>X"00",
4231=>X"00",
4232=>X"00",
4233=>X"00",
4234=>X"00",
4235=>X"00",
4236=>X"00",
4237=>X"00",
4238=>X"00",
4239=>X"00",
4240=>X"00",
4241=>X"00",
4242=>X"00",
4243=>X"00",
4244=>X"00",
4245=>X"00",
4246=>X"00",
4247=>X"00",
4248=>X"00",
4249=>X"00",
4250=>X"00",
4251=>X"00",
4252=>X"00",
4253=>X"00",
4254=>X"00",
4255=>X"00",
4256=>X"00",
4257=>X"00",
4258=>X"00",
4259=>X"00",
4260=>X"00",
4261=>X"00",
4262=>X"00",
4263=>X"00",
4264=>X"00",
4265=>X"00",
4266=>X"00",
4267=>X"00",
4268=>X"00",
4269=>X"00",
4270=>X"00",
4271=>X"00",
4272=>X"00",
4273=>X"00",
4274=>X"00",
4275=>X"00",
4276=>X"00",
4277=>X"00",
4278=>X"00",
4279=>X"00",
4280=>X"00",
4281=>X"00",
4282=>X"00",
4283=>X"00",
4284=>X"00",
4285=>X"00",
4286=>X"00",
4287=>X"00",
4288=>X"00",
4289=>X"00",
4290=>X"00",
4291=>X"00",
4292=>X"00",
4293=>X"00",
4294=>X"00",
4295=>X"00",
4296=>X"00",
4297=>X"00",
4298=>X"00",
4299=>X"00",
4300=>X"00",
4301=>X"00",
4302=>X"00",
4303=>X"00",
4304=>X"00",
4305=>X"00",
4306=>X"00",
4307=>X"00",
4308=>X"00",
4309=>X"00",
4310=>X"00",
4311=>X"00",
4312=>X"00",
4313=>X"00",
4314=>X"00",
4315=>X"00",
4316=>X"00",
4317=>X"00",
4318=>X"00",
4319=>X"00",
4320=>X"00",
4321=>X"00",
4322=>X"00",
4323=>X"00",
4324=>X"00",
4325=>X"00",
4326=>X"00",
4327=>X"00",
4328=>X"00",
4329=>X"00",
4330=>X"00",
4331=>X"00",
4332=>X"00",
4333=>X"00",
4334=>X"00",
4335=>X"00",
4336=>X"00",
4337=>X"00",
4338=>X"00",
4339=>X"00",
4340=>X"00",
4341=>X"00",
4342=>X"00",
4343=>X"00",
4344=>X"00",
4345=>X"00",
4346=>X"00",
4347=>X"00",
4348=>X"00",
4349=>X"00",
4350=>X"00",
4351=>X"00",
4352=>X"15",
4353=>X"15",
4354=>X"15",
4355=>X"15",
4356=>X"15",
4357=>X"15",
4358=>X"15",
4359=>X"15",
4360=>X"15",
4361=>X"15",
4362=>X"15",
4363=>X"15",
4364=>X"15",
4365=>X"15",
4366=>X"15",
4367=>X"15",
4368=>X"15",
4369=>X"15",
4370=>X"15",
4371=>X"15",
4372=>X"15",
4373=>X"15",
4374=>X"15",
4375=>X"15",
4376=>X"15",
4377=>X"15",
4378=>X"15",
4379=>X"15",
4380=>X"19",
4381=>X"19",
4382=>X"15",
4383=>X"15",
4384=>X"15",
4385=>X"15",
4386=>X"19",
4387=>X"19",
4388=>X"15",
4389=>X"15",
4390=>X"15",
4391=>X"15",
4392=>X"19",
4393=>X"19",
4394=>X"15",
4395=>X"15",
4396=>X"19",
4397=>X"19",
4398=>X"25",
4399=>X"25",
4400=>X"29",
4401=>X"29",
4402=>X"3D",
4403=>X"2D",
4404=>X"2D",
4405=>X"29",
4406=>X"2A",
4407=>X"2B",
4408=>X"1B",
4409=>X"1B",
4410=>X"2B",
4411=>X"2A",
4412=>X"25",
4413=>X"34",
4414=>X"34",
4415=>X"35",
4416=>X"35",
4417=>X"25",
4418=>X"25",
4419=>X"25",
4420=>X"25",
4421=>X"25",
4422=>X"25",
4423=>X"25",
4424=>X"25",
4425=>X"25",
4426=>X"25",
4427=>X"25",
4428=>X"25",
4429=>X"25",
4430=>X"15",
4431=>X"15",
4432=>X"15",
4433=>X"15",
4434=>X"15",
4435=>X"15",
4436=>X"15",
4437=>X"15",
4438=>X"15",
4439=>X"15",
4440=>X"15",
4441=>X"15",
4442=>X"15",
4443=>X"15",
4444=>X"15",
4445=>X"15",
4446=>X"15",
4447=>X"15",
4448=>X"15",
4449=>X"15",
4450=>X"15",
4451=>X"15",
4452=>X"00",
4453=>X"00",
4454=>X"00",
4455=>X"00",
4456=>X"00",
4457=>X"00",
4458=>X"00",
4459=>X"00",
4460=>X"00",
4461=>X"00",
4462=>X"00",
4463=>X"00",
4464=>X"00",
4465=>X"00",
4466=>X"00",
4467=>X"00",
4468=>X"00",
4469=>X"00",
4470=>X"00",
4471=>X"00",
4472=>X"00",
4473=>X"00",
4474=>X"00",
4475=>X"00",
4476=>X"00",
4477=>X"00",
4478=>X"00",
4479=>X"00",
4480=>X"00",
4481=>X"00",
4482=>X"00",
4483=>X"00",
4484=>X"00",
4485=>X"00",
4486=>X"00",
4487=>X"00",
4488=>X"00",
4489=>X"00",
4490=>X"00",
4491=>X"00",
4492=>X"00",
4493=>X"00",
4494=>X"00",
4495=>X"00",
4496=>X"00",
4497=>X"00",
4498=>X"00",
4499=>X"00",
4500=>X"00",
4501=>X"00",
4502=>X"00",
4503=>X"00",
4504=>X"00",
4505=>X"00",
4506=>X"00",
4507=>X"00",
4508=>X"00",
4509=>X"00",
4510=>X"00",
4511=>X"00",
4512=>X"00",
4513=>X"00",
4514=>X"00",
4515=>X"00",
4516=>X"00",
4517=>X"00",
4518=>X"00",
4519=>X"00",
4520=>X"00",
4521=>X"00",
4522=>X"00",
4523=>X"00",
4524=>X"00",
4525=>X"00",
4526=>X"00",
4527=>X"00",
4528=>X"00",
4529=>X"00",
4530=>X"00",
4531=>X"00",
4532=>X"00",
4533=>X"00",
4534=>X"00",
4535=>X"00",
4536=>X"00",
4537=>X"00",
4538=>X"00",
4539=>X"00",
4540=>X"00",
4541=>X"00",
4542=>X"00",
4543=>X"00",
4544=>X"00",
4545=>X"00",
4546=>X"00",
4547=>X"00",
4548=>X"00",
4549=>X"00",
4550=>X"00",
4551=>X"00",
4552=>X"00",
4553=>X"00",
4554=>X"00",
4555=>X"00",
4556=>X"00",
4557=>X"00",
4558=>X"00",
4559=>X"00",
4560=>X"00",
4561=>X"00",
4562=>X"00",
4563=>X"00",
4564=>X"00",
4565=>X"00",
4566=>X"00",
4567=>X"00",
4568=>X"00",
4569=>X"00",
4570=>X"00",
4571=>X"00",
4572=>X"00",
4573=>X"00",
4574=>X"00",
4575=>X"00",
4576=>X"00",
4577=>X"00",
4578=>X"00",
4579=>X"00",
4580=>X"00",
4581=>X"00",
4582=>X"00",
4583=>X"00",
4584=>X"00",
4585=>X"00",
4586=>X"00",
4587=>X"00",
4588=>X"00",
4589=>X"00",
4590=>X"00",
4591=>X"00",
4592=>X"00",
4593=>X"00",
4594=>X"00",
4595=>X"00",
4596=>X"00",
4597=>X"00",
4598=>X"00",
4599=>X"00",
4600=>X"00",
4601=>X"00",
4602=>X"00",
4603=>X"00",
4604=>X"00",
4605=>X"00",
4606=>X"00",
4607=>X"00",
4608=>X"15",
4609=>X"15",
4610=>X"15",
4611=>X"15",
4612=>X"15",
4613=>X"15",
4614=>X"15",
4615=>X"15",
4616=>X"15",
4617=>X"15",
4618=>X"15",
4619=>X"15",
4620=>X"15",
4621=>X"15",
4622=>X"15",
4623=>X"15",
4624=>X"15",
4625=>X"15",
4626=>X"15",
4627=>X"15",
4628=>X"15",
4629=>X"15",
4630=>X"15",
4631=>X"15",
4632=>X"15",
4633=>X"15",
4634=>X"19",
4635=>X"15",
4636=>X"15",
4637=>X"19",
4638=>X"15",
4639=>X"19",
4640=>X"15",
4641=>X"19",
4642=>X"15",
4643=>X"19",
4644=>X"15",
4645=>X"19",
4646=>X"15",
4647=>X"19",
4648=>X"15",
4649=>X"19",
4650=>X"15",
4651=>X"19",
4652=>X"15",
4653=>X"19",
4654=>X"25",
4655=>X"29",
4656=>X"2D",
4657=>X"3D",
4658=>X"3C",
4659=>X"2C",
4660=>X"28",
4661=>X"29",
4662=>X"29",
4663=>X"1A",
4664=>X"1B",
4665=>X"1B",
4666=>X"1B",
4667=>X"2A",
4668=>X"25",
4669=>X"25",
4670=>X"35",
4671=>X"35",
4672=>X"35",
4673=>X"39",
4674=>X"26",
4675=>X"25",
4676=>X"25",
4677=>X"25",
4678=>X"25",
4679=>X"25",
4680=>X"15",
4681=>X"25",
4682=>X"15",
4683=>X"25",
4684=>X"15",
4685=>X"25",
4686=>X"15",
4687=>X"15",
4688=>X"25",
4689=>X"15",
4690=>X"15",
4691=>X"15",
4692=>X"25",
4693=>X"15",
4694=>X"15",
4695=>X"25",
4696=>X"15",
4697=>X"15",
4698=>X"15",
4699=>X"15",
4700=>X"15",
4701=>X"15",
4702=>X"15",
4703=>X"15",
4704=>X"15",
4705=>X"15",
4706=>X"15",
4707=>X"15",
4708=>X"00",
4709=>X"00",
4710=>X"00",
4711=>X"00",
4712=>X"00",
4713=>X"00",
4714=>X"00",
4715=>X"00",
4716=>X"00",
4717=>X"00",
4718=>X"00",
4719=>X"00",
4720=>X"00",
4721=>X"00",
4722=>X"00",
4723=>X"00",
4724=>X"00",
4725=>X"00",
4726=>X"00",
4727=>X"00",
4728=>X"00",
4729=>X"00",
4730=>X"00",
4731=>X"00",
4732=>X"00",
4733=>X"00",
4734=>X"00",
4735=>X"00",
4736=>X"00",
4737=>X"00",
4738=>X"00",
4739=>X"00",
4740=>X"00",
4741=>X"00",
4742=>X"00",
4743=>X"00",
4744=>X"00",
4745=>X"00",
4746=>X"00",
4747=>X"00",
4748=>X"00",
4749=>X"00",
4750=>X"00",
4751=>X"00",
4752=>X"00",
4753=>X"00",
4754=>X"00",
4755=>X"00",
4756=>X"00",
4757=>X"00",
4758=>X"00",
4759=>X"00",
4760=>X"00",
4761=>X"00",
4762=>X"00",
4763=>X"00",
4764=>X"00",
4765=>X"00",
4766=>X"00",
4767=>X"00",
4768=>X"00",
4769=>X"00",
4770=>X"00",
4771=>X"00",
4772=>X"00",
4773=>X"00",
4774=>X"00",
4775=>X"00",
4776=>X"00",
4777=>X"00",
4778=>X"00",
4779=>X"00",
4780=>X"00",
4781=>X"00",
4782=>X"00",
4783=>X"00",
4784=>X"00",
4785=>X"00",
4786=>X"00",
4787=>X"00",
4788=>X"00",
4789=>X"00",
4790=>X"00",
4791=>X"00",
4792=>X"00",
4793=>X"00",
4794=>X"00",
4795=>X"00",
4796=>X"00",
4797=>X"00",
4798=>X"00",
4799=>X"00",
4800=>X"00",
4801=>X"00",
4802=>X"00",
4803=>X"00",
4804=>X"00",
4805=>X"00",
4806=>X"00",
4807=>X"00",
4808=>X"00",
4809=>X"00",
4810=>X"00",
4811=>X"00",
4812=>X"00",
4813=>X"00",
4814=>X"00",
4815=>X"00",
4816=>X"00",
4817=>X"00",
4818=>X"00",
4819=>X"00",
4820=>X"00",
4821=>X"00",
4822=>X"00",
4823=>X"00",
4824=>X"00",
4825=>X"00",
4826=>X"00",
4827=>X"00",
4828=>X"00",
4829=>X"00",
4830=>X"00",
4831=>X"00",
4832=>X"00",
4833=>X"00",
4834=>X"00",
4835=>X"00",
4836=>X"00",
4837=>X"00",
4838=>X"00",
4839=>X"00",
4840=>X"00",
4841=>X"00",
4842=>X"00",
4843=>X"00",
4844=>X"00",
4845=>X"00",
4846=>X"00",
4847=>X"00",
4848=>X"00",
4849=>X"00",
4850=>X"00",
4851=>X"00",
4852=>X"00",
4853=>X"00",
4854=>X"00",
4855=>X"00",
4856=>X"00",
4857=>X"00",
4858=>X"00",
4859=>X"00",
4860=>X"00",
4861=>X"00",
4862=>X"00",
4863=>X"00",
4864=>X"15",
4865=>X"15",
4866=>X"15",
4867=>X"15",
4868=>X"15",
4869=>X"15",
4870=>X"15",
4871=>X"15",
4872=>X"15",
4873=>X"15",
4874=>X"15",
4875=>X"15",
4876=>X"15",
4877=>X"15",
4878=>X"15",
4879=>X"15",
4880=>X"15",
4881=>X"15",
4882=>X"15",
4883=>X"15",
4884=>X"15",
4885=>X"15",
4886=>X"15",
4887=>X"15",
4888=>X"15",
4889=>X"15",
4890=>X"15",
4891=>X"15",
4892=>X"19",
4893=>X"15",
4894=>X"15",
4895=>X"15",
4896=>X"15",
4897=>X"15",
4898=>X"15",
4899=>X"15",
4900=>X"19",
4901=>X"19",
4902=>X"15",
4903=>X"15",
4904=>X"15",
4905=>X"15",
4906=>X"19",
4907=>X"19",
4908=>X"15",
4909=>X"15",
4910=>X"29",
4911=>X"3D",
4912=>X"3D",
4913=>X"3C",
4914=>X"28",
4915=>X"29",
4916=>X"29",
4917=>X"19",
4918=>X"19",
4919=>X"19",
4920=>X"1B",
4921=>X"1B",
4922=>X"1B",
4923=>X"26",
4924=>X"35",
4925=>X"25",
4926=>X"25",
4927=>X"25",
4928=>X"35",
4929=>X"3A",
4930=>X"3A",
4931=>X"2A",
4932=>X"29",
4933=>X"25",
4934=>X"25",
4935=>X"25",
4936=>X"25",
4937=>X"25",
4938=>X"15",
4939=>X"25",
4940=>X"15",
4941=>X"25",
4942=>X"15",
4943=>X"15",
4944=>X"15",
4945=>X"15",
4946=>X"15",
4947=>X"15",
4948=>X"15",
4949=>X"15",
4950=>X"15",
4951=>X"15",
4952=>X"15",
4953=>X"15",
4954=>X"15",
4955=>X"15",
4956=>X"15",
4957=>X"15",
4958=>X"15",
4959=>X"15",
4960=>X"15",
4961=>X"15",
4962=>X"15",
4963=>X"15",
4964=>X"00",
4965=>X"00",
4966=>X"00",
4967=>X"00",
4968=>X"00",
4969=>X"00",
4970=>X"00",
4971=>X"00",
4972=>X"00",
4973=>X"00",
4974=>X"00",
4975=>X"00",
4976=>X"00",
4977=>X"00",
4978=>X"00",
4979=>X"00",
4980=>X"00",
4981=>X"00",
4982=>X"00",
4983=>X"00",
4984=>X"00",
4985=>X"00",
4986=>X"00",
4987=>X"00",
4988=>X"00",
4989=>X"00",
4990=>X"00",
4991=>X"00",
4992=>X"00",
4993=>X"00",
4994=>X"00",
4995=>X"00",
4996=>X"00",
4997=>X"00",
4998=>X"00",
4999=>X"00",
5000=>X"00",
5001=>X"00",
5002=>X"00",
5003=>X"00",
5004=>X"00",
5005=>X"00",
5006=>X"00",
5007=>X"00",
5008=>X"00",
5009=>X"00",
5010=>X"00",
5011=>X"00",
5012=>X"00",
5013=>X"00",
5014=>X"00",
5015=>X"00",
5016=>X"00",
5017=>X"00",
5018=>X"00",
5019=>X"00",
5020=>X"00",
5021=>X"00",
5022=>X"00",
5023=>X"00",
5024=>X"00",
5025=>X"00",
5026=>X"00",
5027=>X"00",
5028=>X"00",
5029=>X"00",
5030=>X"00",
5031=>X"00",
5032=>X"00",
5033=>X"00",
5034=>X"00",
5035=>X"00",
5036=>X"00",
5037=>X"00",
5038=>X"00",
5039=>X"00",
5040=>X"00",
5041=>X"00",
5042=>X"00",
5043=>X"00",
5044=>X"00",
5045=>X"00",
5046=>X"00",
5047=>X"00",
5048=>X"00",
5049=>X"00",
5050=>X"00",
5051=>X"00",
5052=>X"00",
5053=>X"00",
5054=>X"00",
5055=>X"00",
5056=>X"00",
5057=>X"00",
5058=>X"00",
5059=>X"00",
5060=>X"00",
5061=>X"00",
5062=>X"00",
5063=>X"00",
5064=>X"00",
5065=>X"00",
5066=>X"00",
5067=>X"00",
5068=>X"00",
5069=>X"00",
5070=>X"00",
5071=>X"00",
5072=>X"00",
5073=>X"00",
5074=>X"00",
5075=>X"00",
5076=>X"00",
5077=>X"00",
5078=>X"00",
5079=>X"00",
5080=>X"00",
5081=>X"00",
5082=>X"00",
5083=>X"00",
5084=>X"00",
5085=>X"00",
5086=>X"00",
5087=>X"00",
5088=>X"00",
5089=>X"00",
5090=>X"00",
5091=>X"00",
5092=>X"00",
5093=>X"00",
5094=>X"00",
5095=>X"00",
5096=>X"00",
5097=>X"00",
5098=>X"00",
5099=>X"00",
5100=>X"00",
5101=>X"00",
5102=>X"00",
5103=>X"00",
5104=>X"00",
5105=>X"00",
5106=>X"00",
5107=>X"00",
5108=>X"00",
5109=>X"00",
5110=>X"00",
5111=>X"00",
5112=>X"00",
5113=>X"00",
5114=>X"00",
5115=>X"00",
5116=>X"00",
5117=>X"00",
5118=>X"00",
5119=>X"00",
5120=>X"15",
5121=>X"15",
5122=>X"15",
5123=>X"15",
5124=>X"15",
5125=>X"15",
5126=>X"15",
5127=>X"15",
5128=>X"15",
5129=>X"15",
5130=>X"15",
5131=>X"15",
5132=>X"15",
5133=>X"15",
5134=>X"15",
5135=>X"15",
5136=>X"15",
5137=>X"15",
5138=>X"15",
5139=>X"15",
5140=>X"15",
5141=>X"15",
5142=>X"15",
5143=>X"15",
5144=>X"15",
5145=>X"15",
5146=>X"15",
5147=>X"15",
5148=>X"19",
5149=>X"15",
5150=>X"19",
5151=>X"15",
5152=>X"19",
5153=>X"15",
5154=>X"15",
5155=>X"15",
5156=>X"19",
5157=>X"15",
5158=>X"19",
5159=>X"15",
5160=>X"19",
5161=>X"15",
5162=>X"19",
5163=>X"15",
5164=>X"15",
5165=>X"29",
5166=>X"29",
5167=>X"3D",
5168=>X"3D",
5169=>X"29",
5170=>X"28",
5171=>X"29",
5172=>X"19",
5173=>X"19",
5174=>X"29",
5175=>X"19",
5176=>X"1B",
5177=>X"1F",
5178=>X"2B",
5179=>X"26",
5180=>X"25",
5181=>X"25",
5182=>X"15",
5183=>X"25",
5184=>X"25",
5185=>X"35",
5186=>X"3F",
5187=>X"3F",
5188=>X"3E",
5189=>X"2A",
5190=>X"29",
5191=>X"25",
5192=>X"25",
5193=>X"25",
5194=>X"15",
5195=>X"25",
5196=>X"15",
5197=>X"25",
5198=>X"15",
5199=>X"15",
5200=>X"15",
5201=>X"15",
5202=>X"15",
5203=>X"25",
5204=>X"15",
5205=>X"15",
5206=>X"15",
5207=>X"15",
5208=>X"15",
5209=>X"15",
5210=>X"15",
5211=>X"15",
5212=>X"15",
5213=>X"15",
5214=>X"15",
5215=>X"15",
5216=>X"15",
5217=>X"15",
5218=>X"15",
5219=>X"15",
5220=>X"00",
5221=>X"00",
5222=>X"00",
5223=>X"00",
5224=>X"00",
5225=>X"00",
5226=>X"00",
5227=>X"00",
5228=>X"00",
5229=>X"00",
5230=>X"00",
5231=>X"00",
5232=>X"00",
5233=>X"00",
5234=>X"00",
5235=>X"00",
5236=>X"00",
5237=>X"00",
5238=>X"00",
5239=>X"00",
5240=>X"00",
5241=>X"00",
5242=>X"00",
5243=>X"00",
5244=>X"00",
5245=>X"00",
5246=>X"00",
5247=>X"00",
5248=>X"00",
5249=>X"00",
5250=>X"00",
5251=>X"00",
5252=>X"00",
5253=>X"00",
5254=>X"00",
5255=>X"00",
5256=>X"00",
5257=>X"00",
5258=>X"00",
5259=>X"00",
5260=>X"00",
5261=>X"00",
5262=>X"00",
5263=>X"00",
5264=>X"00",
5265=>X"00",
5266=>X"00",
5267=>X"00",
5268=>X"00",
5269=>X"00",
5270=>X"00",
5271=>X"00",
5272=>X"00",
5273=>X"00",
5274=>X"00",
5275=>X"00",
5276=>X"00",
5277=>X"00",
5278=>X"00",
5279=>X"00",
5280=>X"00",
5281=>X"00",
5282=>X"00",
5283=>X"00",
5284=>X"00",
5285=>X"00",
5286=>X"00",
5287=>X"00",
5288=>X"00",
5289=>X"00",
5290=>X"00",
5291=>X"00",
5292=>X"00",
5293=>X"00",
5294=>X"00",
5295=>X"00",
5296=>X"00",
5297=>X"00",
5298=>X"00",
5299=>X"00",
5300=>X"00",
5301=>X"00",
5302=>X"00",
5303=>X"00",
5304=>X"00",
5305=>X"00",
5306=>X"00",
5307=>X"00",
5308=>X"00",
5309=>X"00",
5310=>X"00",
5311=>X"00",
5312=>X"00",
5313=>X"00",
5314=>X"00",
5315=>X"00",
5316=>X"00",
5317=>X"00",
5318=>X"00",
5319=>X"00",
5320=>X"00",
5321=>X"00",
5322=>X"00",
5323=>X"00",
5324=>X"00",
5325=>X"00",
5326=>X"00",
5327=>X"00",
5328=>X"00",
5329=>X"00",
5330=>X"00",
5331=>X"00",
5332=>X"00",
5333=>X"00",
5334=>X"00",
5335=>X"00",
5336=>X"00",
5337=>X"00",
5338=>X"00",
5339=>X"00",
5340=>X"00",
5341=>X"00",
5342=>X"00",
5343=>X"00",
5344=>X"00",
5345=>X"00",
5346=>X"00",
5347=>X"00",
5348=>X"00",
5349=>X"00",
5350=>X"00",
5351=>X"00",
5352=>X"00",
5353=>X"00",
5354=>X"00",
5355=>X"00",
5356=>X"00",
5357=>X"00",
5358=>X"00",
5359=>X"00",
5360=>X"00",
5361=>X"00",
5362=>X"00",
5363=>X"00",
5364=>X"00",
5365=>X"00",
5366=>X"00",
5367=>X"00",
5368=>X"00",
5369=>X"00",
5370=>X"00",
5371=>X"00",
5372=>X"00",
5373=>X"00",
5374=>X"00",
5375=>X"00",
5376=>X"15",
5377=>X"15",
5378=>X"15",
5379=>X"15",
5380=>X"15",
5381=>X"15",
5382=>X"15",
5383=>X"15",
5384=>X"15",
5385=>X"15",
5386=>X"15",
5387=>X"15",
5388=>X"15",
5389=>X"15",
5390=>X"15",
5391=>X"15",
5392=>X"15",
5393=>X"15",
5394=>X"15",
5395=>X"15",
5396=>X"15",
5397=>X"15",
5398=>X"15",
5399=>X"19",
5400=>X"15",
5401=>X"15",
5402=>X"15",
5403=>X"15",
5404=>X"15",
5405=>X"15",
5406=>X"19",
5407=>X"15",
5408=>X"19",
5409=>X"15",
5410=>X"15",
5411=>X"19",
5412=>X"15",
5413=>X"15",
5414=>X"19",
5415=>X"15",
5416=>X"19",
5417=>X"15",
5418=>X"19",
5419=>X"15",
5420=>X"29",
5421=>X"29",
5422=>X"29",
5423=>X"29",
5424=>X"29",
5425=>X"29",
5426=>X"29",
5427=>X"19",
5428=>X"19",
5429=>X"19",
5430=>X"29",
5431=>X"19",
5432=>X"1B",
5433=>X"1F",
5434=>X"2B",
5435=>X"26",
5436=>X"25",
5437=>X"25",
5438=>X"25",
5439=>X"15",
5440=>X"25",
5441=>X"25",
5442=>X"3A",
5443=>X"3F",
5444=>X"3F",
5445=>X"3F",
5446=>X"2A",
5447=>X"2A",
5448=>X"25",
5449=>X"25",
5450=>X"15",
5451=>X"25",
5452=>X"25",
5453=>X"15",
5454=>X"15",
5455=>X"15",
5456=>X"15",
5457=>X"15",
5458=>X"15",
5459=>X"25",
5460=>X"15",
5461=>X"15",
5462=>X"15",
5463=>X"15",
5464=>X"15",
5465=>X"15",
5466=>X"15",
5467=>X"15",
5468=>X"15",
5469=>X"15",
5470=>X"15",
5471=>X"15",
5472=>X"15",
5473=>X"15",
5474=>X"15",
5475=>X"15",
5476=>X"00",
5477=>X"00",
5478=>X"00",
5479=>X"00",
5480=>X"00",
5481=>X"00",
5482=>X"00",
5483=>X"00",
5484=>X"00",
5485=>X"00",
5486=>X"00",
5487=>X"00",
5488=>X"00",
5489=>X"00",
5490=>X"00",
5491=>X"00",
5492=>X"00",
5493=>X"00",
5494=>X"00",
5495=>X"00",
5496=>X"00",
5497=>X"00",
5498=>X"00",
5499=>X"00",
5500=>X"00",
5501=>X"00",
5502=>X"00",
5503=>X"00",
5504=>X"00",
5505=>X"00",
5506=>X"00",
5507=>X"00",
5508=>X"00",
5509=>X"00",
5510=>X"00",
5511=>X"00",
5512=>X"00",
5513=>X"00",
5514=>X"00",
5515=>X"00",
5516=>X"00",
5517=>X"00",
5518=>X"00",
5519=>X"00",
5520=>X"00",
5521=>X"00",
5522=>X"00",
5523=>X"00",
5524=>X"00",
5525=>X"00",
5526=>X"00",
5527=>X"00",
5528=>X"00",
5529=>X"00",
5530=>X"00",
5531=>X"00",
5532=>X"00",
5533=>X"00",
5534=>X"00",
5535=>X"00",
5536=>X"00",
5537=>X"00",
5538=>X"00",
5539=>X"00",
5540=>X"00",
5541=>X"00",
5542=>X"00",
5543=>X"00",
5544=>X"00",
5545=>X"00",
5546=>X"00",
5547=>X"00",
5548=>X"00",
5549=>X"00",
5550=>X"00",
5551=>X"00",
5552=>X"00",
5553=>X"00",
5554=>X"00",
5555=>X"00",
5556=>X"00",
5557=>X"00",
5558=>X"00",
5559=>X"00",
5560=>X"00",
5561=>X"00",
5562=>X"00",
5563=>X"00",
5564=>X"00",
5565=>X"00",
5566=>X"00",
5567=>X"00",
5568=>X"00",
5569=>X"00",
5570=>X"00",
5571=>X"00",
5572=>X"00",
5573=>X"00",
5574=>X"00",
5575=>X"00",
5576=>X"00",
5577=>X"00",
5578=>X"00",
5579=>X"00",
5580=>X"00",
5581=>X"00",
5582=>X"00",
5583=>X"00",
5584=>X"00",
5585=>X"00",
5586=>X"00",
5587=>X"00",
5588=>X"00",
5589=>X"00",
5590=>X"00",
5591=>X"00",
5592=>X"00",
5593=>X"00",
5594=>X"00",
5595=>X"00",
5596=>X"00",
5597=>X"00",
5598=>X"00",
5599=>X"00",
5600=>X"00",
5601=>X"00",
5602=>X"00",
5603=>X"00",
5604=>X"00",
5605=>X"00",
5606=>X"00",
5607=>X"00",
5608=>X"00",
5609=>X"00",
5610=>X"00",
5611=>X"00",
5612=>X"00",
5613=>X"00",
5614=>X"00",
5615=>X"00",
5616=>X"00",
5617=>X"00",
5618=>X"00",
5619=>X"00",
5620=>X"00",
5621=>X"00",
5622=>X"00",
5623=>X"00",
5624=>X"00",
5625=>X"00",
5626=>X"00",
5627=>X"00",
5628=>X"00",
5629=>X"00",
5630=>X"00",
5631=>X"00",
5632=>X"15",
5633=>X"15",
5634=>X"15",
5635=>X"15",
5636=>X"15",
5637=>X"15",
5638=>X"15",
5639=>X"15",
5640=>X"15",
5641=>X"15",
5642=>X"15",
5643=>X"15",
5644=>X"15",
5645=>X"15",
5646=>X"15",
5647=>X"15",
5648=>X"15",
5649=>X"15",
5650=>X"15",
5651=>X"15",
5652=>X"15",
5653=>X"15",
5654=>X"19",
5655=>X"19",
5656=>X"15",
5657=>X"19",
5658=>X"15",
5659=>X"19",
5660=>X"15",
5661=>X"15",
5662=>X"19",
5663=>X"15",
5664=>X"19",
5665=>X"15",
5666=>X"15",
5667=>X"19",
5668=>X"15",
5669=>X"15",
5670=>X"19",
5671=>X"15",
5672=>X"19",
5673=>X"15",
5674=>X"19",
5675=>X"29",
5676=>X"29",
5677=>X"29",
5678=>X"29",
5679=>X"29",
5680=>X"29",
5681=>X"29",
5682=>X"19",
5683=>X"19",
5684=>X"19",
5685=>X"19",
5686=>X"19",
5687=>X"19",
5688=>X"1B",
5689=>X"1B",
5690=>X"2A",
5691=>X"25",
5692=>X"25",
5693=>X"25",
5694=>X"25",
5695=>X"25",
5696=>X"25",
5697=>X"25",
5698=>X"2A",
5699=>X"3A",
5700=>X"3F",
5701=>X"3F",
5702=>X"3F",
5703=>X"3A",
5704=>X"25",
5705=>X"25",
5706=>X"15",
5707=>X"25",
5708=>X"25",
5709=>X"15",
5710=>X"15",
5711=>X"15",
5712=>X"15",
5713=>X"15",
5714=>X"15",
5715=>X"15",
5716=>X"15",
5717=>X"15",
5718=>X"15",
5719=>X"15",
5720=>X"15",
5721=>X"15",
5722=>X"15",
5723=>X"15",
5724=>X"15",
5725=>X"15",
5726=>X"15",
5727=>X"15",
5728=>X"15",
5729=>X"15",
5730=>X"15",
5731=>X"15",
5732=>X"00",
5733=>X"00",
5734=>X"00",
5735=>X"00",
5736=>X"00",
5737=>X"00",
5738=>X"00",
5739=>X"00",
5740=>X"00",
5741=>X"00",
5742=>X"00",
5743=>X"00",
5744=>X"00",
5745=>X"00",
5746=>X"00",
5747=>X"00",
5748=>X"00",
5749=>X"00",
5750=>X"00",
5751=>X"00",
5752=>X"00",
5753=>X"00",
5754=>X"00",
5755=>X"00",
5756=>X"00",
5757=>X"00",
5758=>X"00",
5759=>X"00",
5760=>X"00",
5761=>X"00",
5762=>X"00",
5763=>X"00",
5764=>X"00",
5765=>X"00",
5766=>X"00",
5767=>X"00",
5768=>X"00",
5769=>X"00",
5770=>X"00",
5771=>X"00",
5772=>X"00",
5773=>X"00",
5774=>X"00",
5775=>X"00",
5776=>X"00",
5777=>X"00",
5778=>X"00",
5779=>X"00",
5780=>X"00",
5781=>X"00",
5782=>X"00",
5783=>X"00",
5784=>X"00",
5785=>X"00",
5786=>X"00",
5787=>X"00",
5788=>X"00",
5789=>X"00",
5790=>X"00",
5791=>X"00",
5792=>X"00",
5793=>X"00",
5794=>X"00",
5795=>X"00",
5796=>X"00",
5797=>X"00",
5798=>X"00",
5799=>X"00",
5800=>X"00",
5801=>X"00",
5802=>X"00",
5803=>X"00",
5804=>X"00",
5805=>X"00",
5806=>X"00",
5807=>X"00",
5808=>X"00",
5809=>X"00",
5810=>X"00",
5811=>X"00",
5812=>X"00",
5813=>X"00",
5814=>X"00",
5815=>X"00",
5816=>X"00",
5817=>X"00",
5818=>X"00",
5819=>X"00",
5820=>X"00",
5821=>X"00",
5822=>X"00",
5823=>X"00",
5824=>X"00",
5825=>X"00",
5826=>X"00",
5827=>X"00",
5828=>X"00",
5829=>X"00",
5830=>X"00",
5831=>X"00",
5832=>X"00",
5833=>X"00",
5834=>X"00",
5835=>X"00",
5836=>X"00",
5837=>X"00",
5838=>X"00",
5839=>X"00",
5840=>X"00",
5841=>X"00",
5842=>X"00",
5843=>X"00",
5844=>X"00",
5845=>X"00",
5846=>X"00",
5847=>X"00",
5848=>X"00",
5849=>X"00",
5850=>X"00",
5851=>X"00",
5852=>X"00",
5853=>X"00",
5854=>X"00",
5855=>X"00",
5856=>X"00",
5857=>X"00",
5858=>X"00",
5859=>X"00",
5860=>X"00",
5861=>X"00",
5862=>X"00",
5863=>X"00",
5864=>X"00",
5865=>X"00",
5866=>X"00",
5867=>X"00",
5868=>X"00",
5869=>X"00",
5870=>X"00",
5871=>X"00",
5872=>X"00",
5873=>X"00",
5874=>X"00",
5875=>X"00",
5876=>X"00",
5877=>X"00",
5878=>X"00",
5879=>X"00",
5880=>X"00",
5881=>X"00",
5882=>X"00",
5883=>X"00",
5884=>X"00",
5885=>X"00",
5886=>X"00",
5887=>X"00",
5888=>X"15",
5889=>X"15",
5890=>X"15",
5891=>X"15",
5892=>X"15",
5893=>X"15",
5894=>X"15",
5895=>X"15",
5896=>X"15",
5897=>X"15",
5898=>X"15",
5899=>X"15",
5900=>X"15",
5901=>X"15",
5902=>X"15",
5903=>X"15",
5904=>X"15",
5905=>X"15",
5906=>X"19",
5907=>X"15",
5908=>X"15",
5909=>X"19",
5910=>X"19",
5911=>X"15",
5912=>X"15",
5913=>X"19",
5914=>X"15",
5915=>X"15",
5916=>X"15",
5917=>X"15",
5918=>X"19",
5919=>X"15",
5920=>X"19",
5921=>X"15",
5922=>X"15",
5923=>X"15",
5924=>X"15",
5925=>X"15",
5926=>X"19",
5927=>X"15",
5928=>X"19",
5929=>X"15",
5930=>X"29",
5931=>X"2A",
5932=>X"29",
5933=>X"29",
5934=>X"29",
5935=>X"29",
5936=>X"29",
5937=>X"29",
5938=>X"29",
5939=>X"19",
5940=>X"19",
5941=>X"19",
5942=>X"19",
5943=>X"1A",
5944=>X"1B",
5945=>X"1B",
5946=>X"26",
5947=>X"25",
5948=>X"20",
5949=>X"25",
5950=>X"25",
5951=>X"25",
5952=>X"25",
5953=>X"2A",
5954=>X"2A",
5955=>X"2A",
5956=>X"2A",
5957=>X"3A",
5958=>X"3A",
5959=>X"3A",
5960=>X"25",
5961=>X"15",
5962=>X"15",
5963=>X"15",
5964=>X"15",
5965=>X"15",
5966=>X"25",
5967=>X"15",
5968=>X"15",
5969=>X"15",
5970=>X"15",
5971=>X"15",
5972=>X"15",
5973=>X"15",
5974=>X"15",
5975=>X"15",
5976=>X"15",
5977=>X"15",
5978=>X"15",
5979=>X"15",
5980=>X"15",
5981=>X"15",
5982=>X"15",
5983=>X"15",
5984=>X"15",
5985=>X"15",
5986=>X"15",
5987=>X"15",
5988=>X"00",
5989=>X"00",
5990=>X"00",
5991=>X"00",
5992=>X"00",
5993=>X"00",
5994=>X"00",
5995=>X"00",
5996=>X"00",
5997=>X"00",
5998=>X"00",
5999=>X"00",
6000=>X"00",
6001=>X"00",
6002=>X"00",
6003=>X"00",
6004=>X"00",
6005=>X"00",
6006=>X"00",
6007=>X"00",
6008=>X"00",
6009=>X"00",
6010=>X"00",
6011=>X"00",
6012=>X"00",
6013=>X"00",
6014=>X"00",
6015=>X"00",
6016=>X"00",
6017=>X"00",
6018=>X"00",
6019=>X"00",
6020=>X"00",
6021=>X"00",
6022=>X"00",
6023=>X"00",
6024=>X"00",
6025=>X"00",
6026=>X"00",
6027=>X"00",
6028=>X"00",
6029=>X"00",
6030=>X"00",
6031=>X"00",
6032=>X"00",
6033=>X"00",
6034=>X"00",
6035=>X"00",
6036=>X"00",
6037=>X"00",
6038=>X"00",
6039=>X"00",
6040=>X"00",
6041=>X"00",
6042=>X"00",
6043=>X"00",
6044=>X"00",
6045=>X"00",
6046=>X"00",
6047=>X"00",
6048=>X"00",
6049=>X"00",
6050=>X"00",
6051=>X"00",
6052=>X"00",
6053=>X"00",
6054=>X"00",
6055=>X"00",
6056=>X"00",
6057=>X"00",
6058=>X"00",
6059=>X"00",
6060=>X"00",
6061=>X"00",
6062=>X"00",
6063=>X"00",
6064=>X"00",
6065=>X"00",
6066=>X"00",
6067=>X"00",
6068=>X"00",
6069=>X"00",
6070=>X"00",
6071=>X"00",
6072=>X"00",
6073=>X"00",
6074=>X"00",
6075=>X"00",
6076=>X"00",
6077=>X"00",
6078=>X"00",
6079=>X"00",
6080=>X"00",
6081=>X"00",
6082=>X"00",
6083=>X"00",
6084=>X"00",
6085=>X"00",
6086=>X"00",
6087=>X"00",
6088=>X"00",
6089=>X"00",
6090=>X"00",
6091=>X"00",
6092=>X"00",
6093=>X"00",
6094=>X"00",
6095=>X"00",
6096=>X"00",
6097=>X"00",
6098=>X"00",
6099=>X"00",
6100=>X"00",
6101=>X"00",
6102=>X"00",
6103=>X"00",
6104=>X"00",
6105=>X"00",
6106=>X"00",
6107=>X"00",
6108=>X"00",
6109=>X"00",
6110=>X"00",
6111=>X"00",
6112=>X"00",
6113=>X"00",
6114=>X"00",
6115=>X"00",
6116=>X"00",
6117=>X"00",
6118=>X"00",
6119=>X"00",
6120=>X"00",
6121=>X"00",
6122=>X"00",
6123=>X"00",
6124=>X"00",
6125=>X"00",
6126=>X"00",
6127=>X"00",
6128=>X"00",
6129=>X"00",
6130=>X"00",
6131=>X"00",
6132=>X"00",
6133=>X"00",
6134=>X"00",
6135=>X"00",
6136=>X"00",
6137=>X"00",
6138=>X"00",
6139=>X"00",
6140=>X"00",
6141=>X"00",
6142=>X"00",
6143=>X"00",
6144=>X"15",
6145=>X"15",
6146=>X"15",
6147=>X"15",
6148=>X"15",
6149=>X"15",
6150=>X"15",
6151=>X"15",
6152=>X"15",
6153=>X"15",
6154=>X"15",
6155=>X"15",
6156=>X"15",
6157=>X"15",
6158=>X"15",
6159=>X"15",
6160=>X"19",
6161=>X"15",
6162=>X"19",
6163=>X"15",
6164=>X"15",
6165=>X"19",
6166=>X"15",
6167=>X"15",
6168=>X"19",
6169=>X"15",
6170=>X"15",
6171=>X"19",
6172=>X"15",
6173=>X"15",
6174=>X"15",
6175=>X"15",
6176=>X"19",
6177=>X"15",
6178=>X"19",
6179=>X"15",
6180=>X"15",
6181=>X"15",
6182=>X"15",
6183=>X"15",
6184=>X"15",
6185=>X"29",
6186=>X"29",
6187=>X"2A",
6188=>X"29",
6189=>X"29",
6190=>X"29",
6191=>X"29",
6192=>X"29",
6193=>X"19",
6194=>X"2A",
6195=>X"29",
6196=>X"1A",
6197=>X"1A",
6198=>X"1A",
6199=>X"1A",
6200=>X"1B",
6201=>X"1B",
6202=>X"16",
6203=>X"15",
6204=>X"20",
6205=>X"20",
6206=>X"20",
6207=>X"20",
6208=>X"25",
6209=>X"2A",
6210=>X"2A",
6211=>X"2A",
6212=>X"15",
6213=>X"25",
6214=>X"25",
6215=>X"25",
6216=>X"25",
6217=>X"15",
6218=>X"15",
6219=>X"15",
6220=>X"15",
6221=>X"15",
6222=>X"25",
6223=>X"15",
6224=>X"15",
6225=>X"15",
6226=>X"15",
6227=>X"15",
6228=>X"15",
6229=>X"15",
6230=>X"15",
6231=>X"15",
6232=>X"15",
6233=>X"15",
6234=>X"15",
6235=>X"15",
6236=>X"15",
6237=>X"15",
6238=>X"15",
6239=>X"15",
6240=>X"15",
6241=>X"15",
6242=>X"15",
6243=>X"15",
6244=>X"00",
6245=>X"00",
6246=>X"00",
6247=>X"00",
6248=>X"00",
6249=>X"00",
6250=>X"00",
6251=>X"00",
6252=>X"00",
6253=>X"00",
6254=>X"00",
6255=>X"00",
6256=>X"00",
6257=>X"00",
6258=>X"00",
6259=>X"00",
6260=>X"00",
6261=>X"00",
6262=>X"00",
6263=>X"00",
6264=>X"00",
6265=>X"00",
6266=>X"00",
6267=>X"00",
6268=>X"00",
6269=>X"00",
6270=>X"00",
6271=>X"00",
6272=>X"00",
6273=>X"00",
6274=>X"00",
6275=>X"00",
6276=>X"00",
6277=>X"00",
6278=>X"00",
6279=>X"00",
6280=>X"00",
6281=>X"00",
6282=>X"00",
6283=>X"00",
6284=>X"00",
6285=>X"00",
6286=>X"00",
6287=>X"00",
6288=>X"00",
6289=>X"00",
6290=>X"00",
6291=>X"00",
6292=>X"00",
6293=>X"00",
6294=>X"00",
6295=>X"00",
6296=>X"00",
6297=>X"00",
6298=>X"00",
6299=>X"00",
6300=>X"00",
6301=>X"00",
6302=>X"00",
6303=>X"00",
6304=>X"00",
6305=>X"00",
6306=>X"00",
6307=>X"00",
6308=>X"00",
6309=>X"00",
6310=>X"00",
6311=>X"00",
6312=>X"00",
6313=>X"00",
6314=>X"00",
6315=>X"00",
6316=>X"00",
6317=>X"00",
6318=>X"00",
6319=>X"00",
6320=>X"00",
6321=>X"00",
6322=>X"00",
6323=>X"00",
6324=>X"00",
6325=>X"00",
6326=>X"00",
6327=>X"00",
6328=>X"00",
6329=>X"00",
6330=>X"00",
6331=>X"00",
6332=>X"00",
6333=>X"00",
6334=>X"00",
6335=>X"00",
6336=>X"00",
6337=>X"00",
6338=>X"00",
6339=>X"00",
6340=>X"00",
6341=>X"00",
6342=>X"00",
6343=>X"00",
6344=>X"00",
6345=>X"00",
6346=>X"00",
6347=>X"00",
6348=>X"00",
6349=>X"00",
6350=>X"00",
6351=>X"00",
6352=>X"00",
6353=>X"00",
6354=>X"00",
6355=>X"00",
6356=>X"00",
6357=>X"00",
6358=>X"00",
6359=>X"00",
6360=>X"00",
6361=>X"00",
6362=>X"00",
6363=>X"00",
6364=>X"00",
6365=>X"00",
6366=>X"00",
6367=>X"00",
6368=>X"00",
6369=>X"00",
6370=>X"00",
6371=>X"00",
6372=>X"00",
6373=>X"00",
6374=>X"00",
6375=>X"00",
6376=>X"00",
6377=>X"00",
6378=>X"00",
6379=>X"00",
6380=>X"00",
6381=>X"00",
6382=>X"00",
6383=>X"00",
6384=>X"00",
6385=>X"00",
6386=>X"00",
6387=>X"00",
6388=>X"00",
6389=>X"00",
6390=>X"00",
6391=>X"00",
6392=>X"00",
6393=>X"00",
6394=>X"00",
6395=>X"00",
6396=>X"00",
6397=>X"00",
6398=>X"00",
6399=>X"00",
6400=>X"15",
6401=>X"15",
6402=>X"15",
6403=>X"15",
6404=>X"15",
6405=>X"15",
6406=>X"15",
6407=>X"15",
6408=>X"15",
6409=>X"15",
6410=>X"15",
6411=>X"14",
6412=>X"15",
6413=>X"15",
6414=>X"15",
6415=>X"15",
6416=>X"19",
6417=>X"15",
6418=>X"15",
6419=>X"15",
6420=>X"15",
6421=>X"15",
6422=>X"15",
6423=>X"15",
6424=>X"19",
6425=>X"15",
6426=>X"15",
6427=>X"19",
6428=>X"15",
6429=>X"15",
6430=>X"15",
6431=>X"15",
6432=>X"15",
6433=>X"15",
6434=>X"19",
6435=>X"15",
6436=>X"15",
6437=>X"15",
6438=>X"15",
6439=>X"15",
6440=>X"29",
6441=>X"29",
6442=>X"29",
6443=>X"29",
6444=>X"29",
6445=>X"29",
6446=>X"29",
6447=>X"19",
6448=>X"29",
6449=>X"29",
6450=>X"2A",
6451=>X"29",
6452=>X"1A",
6453=>X"1A",
6454=>X"1A",
6455=>X"1A",
6456=>X"1B",
6457=>X"1F",
6458=>X"1A",
6459=>X"15",
6460=>X"10",
6461=>X"10",
6462=>X"24",
6463=>X"24",
6464=>X"25",
6465=>X"25",
6466=>X"15",
6467=>X"15",
6468=>X"15",
6469=>X"15",
6470=>X"15",
6471=>X"15",
6472=>X"15",
6473=>X"15",
6474=>X"15",
6475=>X"15",
6476=>X"15",
6477=>X"15",
6478=>X"15",
6479=>X"15",
6480=>X"15",
6481=>X"15",
6482=>X"15",
6483=>X"15",
6484=>X"15",
6485=>X"15",
6486=>X"15",
6487=>X"15",
6488=>X"15",
6489=>X"15",
6490=>X"15",
6491=>X"15",
6492=>X"15",
6493=>X"15",
6494=>X"15",
6495=>X"15",
6496=>X"15",
6497=>X"15",
6498=>X"15",
6499=>X"15",
6500=>X"00",
6501=>X"00",
6502=>X"00",
6503=>X"00",
6504=>X"00",
6505=>X"00",
6506=>X"00",
6507=>X"00",
6508=>X"00",
6509=>X"00",
6510=>X"00",
6511=>X"00",
6512=>X"00",
6513=>X"00",
6514=>X"00",
6515=>X"00",
6516=>X"00",
6517=>X"00",
6518=>X"00",
6519=>X"00",
6520=>X"00",
6521=>X"00",
6522=>X"00",
6523=>X"00",
6524=>X"00",
6525=>X"00",
6526=>X"00",
6527=>X"00",
6528=>X"00",
6529=>X"00",
6530=>X"00",
6531=>X"00",
6532=>X"00",
6533=>X"00",
6534=>X"00",
6535=>X"00",
6536=>X"00",
6537=>X"00",
6538=>X"00",
6539=>X"00",
6540=>X"00",
6541=>X"00",
6542=>X"00",
6543=>X"00",
6544=>X"00",
6545=>X"00",
6546=>X"00",
6547=>X"00",
6548=>X"00",
6549=>X"00",
6550=>X"00",
6551=>X"00",
6552=>X"00",
6553=>X"00",
6554=>X"00",
6555=>X"00",
6556=>X"00",
6557=>X"00",
6558=>X"00",
6559=>X"00",
6560=>X"00",
6561=>X"00",
6562=>X"00",
6563=>X"00",
6564=>X"00",
6565=>X"00",
6566=>X"00",
6567=>X"00",
6568=>X"00",
6569=>X"00",
6570=>X"00",
6571=>X"00",
6572=>X"00",
6573=>X"00",
6574=>X"00",
6575=>X"00",
6576=>X"00",
6577=>X"00",
6578=>X"00",
6579=>X"00",
6580=>X"00",
6581=>X"00",
6582=>X"00",
6583=>X"00",
6584=>X"00",
6585=>X"00",
6586=>X"00",
6587=>X"00",
6588=>X"00",
6589=>X"00",
6590=>X"00",
6591=>X"00",
6592=>X"00",
6593=>X"00",
6594=>X"00",
6595=>X"00",
6596=>X"00",
6597=>X"00",
6598=>X"00",
6599=>X"00",
6600=>X"00",
6601=>X"00",
6602=>X"00",
6603=>X"00",
6604=>X"00",
6605=>X"00",
6606=>X"00",
6607=>X"00",
6608=>X"00",
6609=>X"00",
6610=>X"00",
6611=>X"00",
6612=>X"00",
6613=>X"00",
6614=>X"00",
6615=>X"00",
6616=>X"00",
6617=>X"00",
6618=>X"00",
6619=>X"00",
6620=>X"00",
6621=>X"00",
6622=>X"00",
6623=>X"00",
6624=>X"00",
6625=>X"00",
6626=>X"00",
6627=>X"00",
6628=>X"00",
6629=>X"00",
6630=>X"00",
6631=>X"00",
6632=>X"00",
6633=>X"00",
6634=>X"00",
6635=>X"00",
6636=>X"00",
6637=>X"00",
6638=>X"00",
6639=>X"00",
6640=>X"00",
6641=>X"00",
6642=>X"00",
6643=>X"00",
6644=>X"00",
6645=>X"00",
6646=>X"00",
6647=>X"00",
6648=>X"00",
6649=>X"00",
6650=>X"00",
6651=>X"00",
6652=>X"00",
6653=>X"00",
6654=>X"00",
6655=>X"00",
6656=>X"15",
6657=>X"15",
6658=>X"15",
6659=>X"15",
6660=>X"15",
6661=>X"15",
6662=>X"15",
6663=>X"15",
6664=>X"15",
6665=>X"15",
6666=>X"14",
6667=>X"14",
6668=>X"15",
6669=>X"15",
6670=>X"15",
6671=>X"15",
6672=>X"15",
6673=>X"15",
6674=>X"15",
6675=>X"15",
6676=>X"15",
6677=>X"15",
6678=>X"19",
6679=>X"15",
6680=>X"15",
6681=>X"15",
6682=>X"15",
6683=>X"15",
6684=>X"15",
6685=>X"19",
6686=>X"15",
6687=>X"15",
6688=>X"15",
6689=>X"15",
6690=>X"15",
6691=>X"15",
6692=>X"15",
6693=>X"15",
6694=>X"19",
6695=>X"29",
6696=>X"2E",
6697=>X"29",
6698=>X"19",
6699=>X"29",
6700=>X"29",
6701=>X"29",
6702=>X"29",
6703=>X"29",
6704=>X"19",
6705=>X"29",
6706=>X"19",
6707=>X"19",
6708=>X"19",
6709=>X"1A",
6710=>X"1A",
6711=>X"1A",
6712=>X"1B",
6713=>X"1B",
6714=>X"1B",
6715=>X"16",
6716=>X"11",
6717=>X"20",
6718=>X"24",
6719=>X"24",
6720=>X"15",
6721=>X"15",
6722=>X"25",
6723=>X"15",
6724=>X"25",
6725=>X"15",
6726=>X"15",
6727=>X"15",
6728=>X"15",
6729=>X"15",
6730=>X"15",
6731=>X"15",
6732=>X"15",
6733=>X"15",
6734=>X"15",
6735=>X"15",
6736=>X"15",
6737=>X"15",
6738=>X"15",
6739=>X"15",
6740=>X"15",
6741=>X"15",
6742=>X"15",
6743=>X"15",
6744=>X"15",
6745=>X"15",
6746=>X"15",
6747=>X"15",
6748=>X"15",
6749=>X"15",
6750=>X"15",
6751=>X"15",
6752=>X"15",
6753=>X"15",
6754=>X"15",
6755=>X"15",
6756=>X"00",
6757=>X"00",
6758=>X"00",
6759=>X"00",
6760=>X"00",
6761=>X"00",
6762=>X"00",
6763=>X"00",
6764=>X"00",
6765=>X"00",
6766=>X"00",
6767=>X"00",
6768=>X"00",
6769=>X"00",
6770=>X"00",
6771=>X"00",
6772=>X"00",
6773=>X"00",
6774=>X"00",
6775=>X"00",
6776=>X"00",
6777=>X"00",
6778=>X"00",
6779=>X"00",
6780=>X"00",
6781=>X"00",
6782=>X"00",
6783=>X"00",
6784=>X"00",
6785=>X"00",
6786=>X"00",
6787=>X"00",
6788=>X"00",
6789=>X"00",
6790=>X"00",
6791=>X"00",
6792=>X"00",
6793=>X"00",
6794=>X"00",
6795=>X"00",
6796=>X"00",
6797=>X"00",
6798=>X"00",
6799=>X"00",
6800=>X"00",
6801=>X"00",
6802=>X"00",
6803=>X"00",
6804=>X"00",
6805=>X"00",
6806=>X"00",
6807=>X"00",
6808=>X"00",
6809=>X"00",
6810=>X"00",
6811=>X"00",
6812=>X"00",
6813=>X"00",
6814=>X"00",
6815=>X"00",
6816=>X"00",
6817=>X"00",
6818=>X"00",
6819=>X"00",
6820=>X"00",
6821=>X"00",
6822=>X"00",
6823=>X"00",
6824=>X"00",
6825=>X"00",
6826=>X"00",
6827=>X"00",
6828=>X"00",
6829=>X"00",
6830=>X"00",
6831=>X"00",
6832=>X"00",
6833=>X"00",
6834=>X"00",
6835=>X"00",
6836=>X"00",
6837=>X"00",
6838=>X"00",
6839=>X"00",
6840=>X"00",
6841=>X"00",
6842=>X"00",
6843=>X"00",
6844=>X"00",
6845=>X"00",
6846=>X"00",
6847=>X"00",
6848=>X"00",
6849=>X"00",
6850=>X"00",
6851=>X"00",
6852=>X"00",
6853=>X"00",
6854=>X"00",
6855=>X"00",
6856=>X"00",
6857=>X"00",
6858=>X"00",
6859=>X"00",
6860=>X"00",
6861=>X"00",
6862=>X"00",
6863=>X"00",
6864=>X"00",
6865=>X"00",
6866=>X"00",
6867=>X"00",
6868=>X"00",
6869=>X"00",
6870=>X"00",
6871=>X"00",
6872=>X"00",
6873=>X"00",
6874=>X"00",
6875=>X"00",
6876=>X"00",
6877=>X"00",
6878=>X"00",
6879=>X"00",
6880=>X"00",
6881=>X"00",
6882=>X"00",
6883=>X"00",
6884=>X"00",
6885=>X"00",
6886=>X"00",
6887=>X"00",
6888=>X"00",
6889=>X"00",
6890=>X"00",
6891=>X"00",
6892=>X"00",
6893=>X"00",
6894=>X"00",
6895=>X"00",
6896=>X"00",
6897=>X"00",
6898=>X"00",
6899=>X"00",
6900=>X"00",
6901=>X"00",
6902=>X"00",
6903=>X"00",
6904=>X"00",
6905=>X"00",
6906=>X"00",
6907=>X"00",
6908=>X"00",
6909=>X"00",
6910=>X"00",
6911=>X"00",
6912=>X"15",
6913=>X"15",
6914=>X"15",
6915=>X"15",
6916=>X"15",
6917=>X"15",
6918=>X"15",
6919=>X"15",
6920=>X"15",
6921=>X"15",
6922=>X"14",
6923=>X"14",
6924=>X"15",
6925=>X"15",
6926=>X"15",
6927=>X"14",
6928=>X"14",
6929=>X"14",
6930=>X"15",
6931=>X"15",
6932=>X"14",
6933=>X"15",
6934=>X"19",
6935=>X"19",
6936=>X"15",
6937=>X"15",
6938=>X"15",
6939=>X"15",
6940=>X"15",
6941=>X"15",
6942=>X"15",
6943=>X"15",
6944=>X"15",
6945=>X"15",
6946=>X"15",
6947=>X"15",
6948=>X"15",
6949=>X"19",
6950=>X"29",
6951=>X"29",
6952=>X"29",
6953=>X"29",
6954=>X"29",
6955=>X"29",
6956=>X"19",
6957=>X"19",
6958=>X"29",
6959=>X"29",
6960=>X"19",
6961=>X"19",
6962=>X"19",
6963=>X"19",
6964=>X"19",
6965=>X"19",
6966=>X"1A",
6967=>X"1A",
6968=>X"1A",
6969=>X"1A",
6970=>X"1B",
6971=>X"1A",
6972=>X"15",
6973=>X"24",
6974=>X"25",
6975=>X"25",
6976=>X"15",
6977=>X"15",
6978=>X"25",
6979=>X"25",
6980=>X"15",
6981=>X"15",
6982=>X"15",
6983=>X"15",
6984=>X"15",
6985=>X"15",
6986=>X"15",
6987=>X"15",
6988=>X"15",
6989=>X"15",
6990=>X"15",
6991=>X"15",
6992=>X"15",
6993=>X"15",
6994=>X"15",
6995=>X"15",
6996=>X"15",
6997=>X"15",
6998=>X"15",
6999=>X"15",
7000=>X"15",
7001=>X"15",
7002=>X"15",
7003=>X"15",
7004=>X"15",
7005=>X"15",
7006=>X"15",
7007=>X"15",
7008=>X"15",
7009=>X"15",
7010=>X"15",
7011=>X"15",
7012=>X"00",
7013=>X"00",
7014=>X"00",
7015=>X"00",
7016=>X"00",
7017=>X"00",
7018=>X"00",
7019=>X"00",
7020=>X"00",
7021=>X"00",
7022=>X"00",
7023=>X"00",
7024=>X"00",
7025=>X"00",
7026=>X"00",
7027=>X"00",
7028=>X"00",
7029=>X"00",
7030=>X"00",
7031=>X"00",
7032=>X"00",
7033=>X"00",
7034=>X"00",
7035=>X"00",
7036=>X"00",
7037=>X"00",
7038=>X"00",
7039=>X"00",
7040=>X"00",
7041=>X"00",
7042=>X"00",
7043=>X"00",
7044=>X"00",
7045=>X"00",
7046=>X"00",
7047=>X"00",
7048=>X"00",
7049=>X"00",
7050=>X"00",
7051=>X"00",
7052=>X"00",
7053=>X"00",
7054=>X"00",
7055=>X"00",
7056=>X"00",
7057=>X"00",
7058=>X"00",
7059=>X"00",
7060=>X"00",
7061=>X"00",
7062=>X"00",
7063=>X"00",
7064=>X"00",
7065=>X"00",
7066=>X"00",
7067=>X"00",
7068=>X"00",
7069=>X"00",
7070=>X"00",
7071=>X"00",
7072=>X"00",
7073=>X"00",
7074=>X"00",
7075=>X"00",
7076=>X"00",
7077=>X"00",
7078=>X"00",
7079=>X"00",
7080=>X"00",
7081=>X"00",
7082=>X"00",
7083=>X"00",
7084=>X"00",
7085=>X"00",
7086=>X"00",
7087=>X"00",
7088=>X"00",
7089=>X"00",
7090=>X"00",
7091=>X"00",
7092=>X"00",
7093=>X"00",
7094=>X"00",
7095=>X"00",
7096=>X"00",
7097=>X"00",
7098=>X"00",
7099=>X"00",
7100=>X"00",
7101=>X"00",
7102=>X"00",
7103=>X"00",
7104=>X"00",
7105=>X"00",
7106=>X"00",
7107=>X"00",
7108=>X"00",
7109=>X"00",
7110=>X"00",
7111=>X"00",
7112=>X"00",
7113=>X"00",
7114=>X"00",
7115=>X"00",
7116=>X"00",
7117=>X"00",
7118=>X"00",
7119=>X"00",
7120=>X"00",
7121=>X"00",
7122=>X"00",
7123=>X"00",
7124=>X"00",
7125=>X"00",
7126=>X"00",
7127=>X"00",
7128=>X"00",
7129=>X"00",
7130=>X"00",
7131=>X"00",
7132=>X"00",
7133=>X"00",
7134=>X"00",
7135=>X"00",
7136=>X"00",
7137=>X"00",
7138=>X"00",
7139=>X"00",
7140=>X"00",
7141=>X"00",
7142=>X"00",
7143=>X"00",
7144=>X"00",
7145=>X"00",
7146=>X"00",
7147=>X"00",
7148=>X"00",
7149=>X"00",
7150=>X"00",
7151=>X"00",
7152=>X"00",
7153=>X"00",
7154=>X"00",
7155=>X"00",
7156=>X"00",
7157=>X"00",
7158=>X"00",
7159=>X"00",
7160=>X"00",
7161=>X"00",
7162=>X"00",
7163=>X"00",
7164=>X"00",
7165=>X"00",
7166=>X"00",
7167=>X"00",
7168=>X"15",
7169=>X"15",
7170=>X"15",
7171=>X"15",
7172=>X"15",
7173=>X"15",
7174=>X"15",
7175=>X"15",
7176=>X"15",
7177=>X"14",
7178=>X"14",
7179=>X"14",
7180=>X"15",
7181=>X"15",
7182=>X"15",
7183=>X"14",
7184=>X"14",
7185=>X"14",
7186=>X"14",
7187=>X"14",
7188=>X"14",
7189=>X"15",
7190=>X"15",
7191=>X"15",
7192=>X"15",
7193=>X"19",
7194=>X"15",
7195=>X"15",
7196=>X"15",
7197=>X"15",
7198=>X"15",
7199=>X"15",
7200=>X"15",
7201=>X"15",
7202=>X"15",
7203=>X"15",
7204=>X"19",
7205=>X"19",
7206=>X"2A",
7207=>X"29",
7208=>X"29",
7209=>X"29",
7210=>X"29",
7211=>X"19",
7212=>X"19",
7213=>X"19",
7214=>X"19",
7215=>X"19",
7216=>X"19",
7217=>X"19",
7218=>X"19",
7219=>X"19",
7220=>X"29",
7221=>X"19",
7222=>X"19",
7223=>X"1A",
7224=>X"1A",
7225=>X"1A",
7226=>X"16",
7227=>X"1B",
7228=>X"16",
7229=>X"16",
7230=>X"25",
7231=>X"15",
7232=>X"15",
7233=>X"19",
7234=>X"15",
7235=>X"15",
7236=>X"15",
7237=>X"15",
7238=>X"15",
7239=>X"15",
7240=>X"15",
7241=>X"15",
7242=>X"15",
7243=>X"15",
7244=>X"15",
7245=>X"25",
7246=>X"15",
7247=>X"15",
7248=>X"15",
7249=>X"15",
7250=>X"15",
7251=>X"15",
7252=>X"15",
7253=>X"15",
7254=>X"15",
7255=>X"15",
7256=>X"15",
7257=>X"15",
7258=>X"15",
7259=>X"15",
7260=>X"15",
7261=>X"15",
7262=>X"15",
7263=>X"15",
7264=>X"15",
7265=>X"15",
7266=>X"15",
7267=>X"15",
7268=>X"00",
7269=>X"00",
7270=>X"00",
7271=>X"00",
7272=>X"00",
7273=>X"00",
7274=>X"00",
7275=>X"00",
7276=>X"00",
7277=>X"00",
7278=>X"00",
7279=>X"00",
7280=>X"00",
7281=>X"00",
7282=>X"00",
7283=>X"00",
7284=>X"00",
7285=>X"00",
7286=>X"00",
7287=>X"00",
7288=>X"00",
7289=>X"00",
7290=>X"00",
7291=>X"00",
7292=>X"00",
7293=>X"00",
7294=>X"00",
7295=>X"00",
7296=>X"00",
7297=>X"00",
7298=>X"00",
7299=>X"00",
7300=>X"00",
7301=>X"00",
7302=>X"00",
7303=>X"00",
7304=>X"00",
7305=>X"00",
7306=>X"00",
7307=>X"00",
7308=>X"00",
7309=>X"00",
7310=>X"00",
7311=>X"00",
7312=>X"00",
7313=>X"00",
7314=>X"00",
7315=>X"00",
7316=>X"00",
7317=>X"00",
7318=>X"00",
7319=>X"00",
7320=>X"00",
7321=>X"00",
7322=>X"00",
7323=>X"00",
7324=>X"00",
7325=>X"00",
7326=>X"00",
7327=>X"00",
7328=>X"00",
7329=>X"00",
7330=>X"00",
7331=>X"00",
7332=>X"00",
7333=>X"00",
7334=>X"00",
7335=>X"00",
7336=>X"00",
7337=>X"00",
7338=>X"00",
7339=>X"00",
7340=>X"00",
7341=>X"00",
7342=>X"00",
7343=>X"00",
7344=>X"00",
7345=>X"00",
7346=>X"00",
7347=>X"00",
7348=>X"00",
7349=>X"00",
7350=>X"00",
7351=>X"00",
7352=>X"00",
7353=>X"00",
7354=>X"00",
7355=>X"00",
7356=>X"00",
7357=>X"00",
7358=>X"00",
7359=>X"00",
7360=>X"00",
7361=>X"00",
7362=>X"00",
7363=>X"00",
7364=>X"00",
7365=>X"00",
7366=>X"00",
7367=>X"00",
7368=>X"00",
7369=>X"00",
7370=>X"00",
7371=>X"00",
7372=>X"00",
7373=>X"00",
7374=>X"00",
7375=>X"00",
7376=>X"00",
7377=>X"00",
7378=>X"00",
7379=>X"00",
7380=>X"00",
7381=>X"00",
7382=>X"00",
7383=>X"00",
7384=>X"00",
7385=>X"00",
7386=>X"00",
7387=>X"00",
7388=>X"00",
7389=>X"00",
7390=>X"00",
7391=>X"00",
7392=>X"00",
7393=>X"00",
7394=>X"00",
7395=>X"00",
7396=>X"00",
7397=>X"00",
7398=>X"00",
7399=>X"00",
7400=>X"00",
7401=>X"00",
7402=>X"00",
7403=>X"00",
7404=>X"00",
7405=>X"00",
7406=>X"00",
7407=>X"00",
7408=>X"00",
7409=>X"00",
7410=>X"00",
7411=>X"00",
7412=>X"00",
7413=>X"00",
7414=>X"00",
7415=>X"00",
7416=>X"00",
7417=>X"00",
7418=>X"00",
7419=>X"00",
7420=>X"00",
7421=>X"00",
7422=>X"00",
7423=>X"00",
7424=>X"15",
7425=>X"15",
7426=>X"15",
7427=>X"15",
7428=>X"15",
7429=>X"15",
7430=>X"15",
7431=>X"15",
7432=>X"15",
7433=>X"14",
7434=>X"14",
7435=>X"14",
7436=>X"14",
7437=>X"14",
7438=>X"14",
7439=>X"14",
7440=>X"14",
7441=>X"14",
7442=>X"14",
7443=>X"14",
7444=>X"14",
7445=>X"15",
7446=>X"15",
7447=>X"15",
7448=>X"15",
7449=>X"15",
7450=>X"15",
7451=>X"15",
7452=>X"19",
7453=>X"15",
7454=>X"15",
7455=>X"15",
7456=>X"15",
7457=>X"15",
7458=>X"15",
7459=>X"15",
7460=>X"19",
7461=>X"2D",
7462=>X"29",
7463=>X"29",
7464=>X"29",
7465=>X"29",
7466=>X"19",
7467=>X"19",
7468=>X"19",
7469=>X"29",
7470=>X"19",
7471=>X"19",
7472=>X"29",
7473=>X"19",
7474=>X"29",
7475=>X"19",
7476=>X"19",
7477=>X"19",
7478=>X"19",
7479=>X"1A",
7480=>X"1A",
7481=>X"1A",
7482=>X"26",
7483=>X"16",
7484=>X"27",
7485=>X"17",
7486=>X"17",
7487=>X"15",
7488=>X"15",
7489=>X"15",
7490=>X"15",
7491=>X"15",
7492=>X"15",
7493=>X"15",
7494=>X"15",
7495=>X"15",
7496=>X"15",
7497=>X"15",
7498=>X"15",
7499=>X"15",
7500=>X"15",
7501=>X"15",
7502=>X"15",
7503=>X"15",
7504=>X"15",
7505=>X"15",
7506=>X"15",
7507=>X"15",
7508=>X"15",
7509=>X"15",
7510=>X"15",
7511=>X"15",
7512=>X"15",
7513=>X"15",
7514=>X"15",
7515=>X"15",
7516=>X"15",
7517=>X"15",
7518=>X"15",
7519=>X"15",
7520=>X"15",
7521=>X"15",
7522=>X"15",
7523=>X"15",
7524=>X"00",
7525=>X"00",
7526=>X"00",
7527=>X"00",
7528=>X"00",
7529=>X"00",
7530=>X"00",
7531=>X"00",
7532=>X"00",
7533=>X"00",
7534=>X"00",
7535=>X"00",
7536=>X"00",
7537=>X"00",
7538=>X"00",
7539=>X"00",
7540=>X"00",
7541=>X"00",
7542=>X"00",
7543=>X"00",
7544=>X"00",
7545=>X"00",
7546=>X"00",
7547=>X"00",
7548=>X"00",
7549=>X"00",
7550=>X"00",
7551=>X"00",
7552=>X"00",
7553=>X"00",
7554=>X"00",
7555=>X"00",
7556=>X"00",
7557=>X"00",
7558=>X"00",
7559=>X"00",
7560=>X"00",
7561=>X"00",
7562=>X"00",
7563=>X"00",
7564=>X"00",
7565=>X"00",
7566=>X"00",
7567=>X"00",
7568=>X"00",
7569=>X"00",
7570=>X"00",
7571=>X"00",
7572=>X"00",
7573=>X"00",
7574=>X"00",
7575=>X"00",
7576=>X"00",
7577=>X"00",
7578=>X"00",
7579=>X"00",
7580=>X"00",
7581=>X"00",
7582=>X"00",
7583=>X"00",
7584=>X"00",
7585=>X"00",
7586=>X"00",
7587=>X"00",
7588=>X"00",
7589=>X"00",
7590=>X"00",
7591=>X"00",
7592=>X"00",
7593=>X"00",
7594=>X"00",
7595=>X"00",
7596=>X"00",
7597=>X"00",
7598=>X"00",
7599=>X"00",
7600=>X"00",
7601=>X"00",
7602=>X"00",
7603=>X"00",
7604=>X"00",
7605=>X"00",
7606=>X"00",
7607=>X"00",
7608=>X"00",
7609=>X"00",
7610=>X"00",
7611=>X"00",
7612=>X"00",
7613=>X"00",
7614=>X"00",
7615=>X"00",
7616=>X"00",
7617=>X"00",
7618=>X"00",
7619=>X"00",
7620=>X"00",
7621=>X"00",
7622=>X"00",
7623=>X"00",
7624=>X"00",
7625=>X"00",
7626=>X"00",
7627=>X"00",
7628=>X"00",
7629=>X"00",
7630=>X"00",
7631=>X"00",
7632=>X"00",
7633=>X"00",
7634=>X"00",
7635=>X"00",
7636=>X"00",
7637=>X"00",
7638=>X"00",
7639=>X"00",
7640=>X"00",
7641=>X"00",
7642=>X"00",
7643=>X"00",
7644=>X"00",
7645=>X"00",
7646=>X"00",
7647=>X"00",
7648=>X"00",
7649=>X"00",
7650=>X"00",
7651=>X"00",
7652=>X"00",
7653=>X"00",
7654=>X"00",
7655=>X"00",
7656=>X"00",
7657=>X"00",
7658=>X"00",
7659=>X"00",
7660=>X"00",
7661=>X"00",
7662=>X"00",
7663=>X"00",
7664=>X"00",
7665=>X"00",
7666=>X"00",
7667=>X"00",
7668=>X"00",
7669=>X"00",
7670=>X"00",
7671=>X"00",
7672=>X"00",
7673=>X"00",
7674=>X"00",
7675=>X"00",
7676=>X"00",
7677=>X"00",
7678=>X"00",
7679=>X"00",
7680=>X"15",
7681=>X"15",
7682=>X"15",
7683=>X"15",
7684=>X"15",
7685=>X"15",
7686=>X"15",
7687=>X"14",
7688=>X"14",
7689=>X"14",
7690=>X"14",
7691=>X"14",
7692=>X"14",
7693=>X"14",
7694=>X"14",
7695=>X"14",
7696=>X"14",
7697=>X"14",
7698=>X"14",
7699=>X"14",
7700=>X"14",
7701=>X"15",
7702=>X"15",
7703=>X"19",
7704=>X"15",
7705=>X"15",
7706=>X"15",
7707=>X"15",
7708=>X"15",
7709=>X"15",
7710=>X"15",
7711=>X"19",
7712=>X"15",
7713=>X"15",
7714=>X"19",
7715=>X"19",
7716=>X"29",
7717=>X"29",
7718=>X"29",
7719=>X"19",
7720=>X"29",
7721=>X"19",
7722=>X"19",
7723=>X"19",
7724=>X"19",
7725=>X"19",
7726=>X"19",
7727=>X"19",
7728=>X"19",
7729=>X"19",
7730=>X"19",
7731=>X"19",
7732=>X"19",
7733=>X"1A",
7734=>X"2A",
7735=>X"1A",
7736=>X"1A",
7737=>X"1A",
7738=>X"1A",
7739=>X"1A",
7740=>X"26",
7741=>X"27",
7742=>X"27",
7743=>X"27",
7744=>X"15",
7745=>X"15",
7746=>X"15",
7747=>X"15",
7748=>X"15",
7749=>X"15",
7750=>X"15",
7751=>X"15",
7752=>X"15",
7753=>X"15",
7754=>X"15",
7755=>X"15",
7756=>X"15",
7757=>X"15",
7758=>X"15",
7759=>X"15",
7760=>X"15",
7761=>X"15",
7762=>X"15",
7763=>X"15",
7764=>X"15",
7765=>X"15",
7766=>X"15",
7767=>X"15",
7768=>X"15",
7769=>X"15",
7770=>X"15",
7771=>X"15",
7772=>X"15",
7773=>X"15",
7774=>X"15",
7775=>X"15",
7776=>X"15",
7777=>X"15",
7778=>X"15",
7779=>X"15",
7780=>X"00",
7781=>X"00",
7782=>X"00",
7783=>X"00",
7784=>X"00",
7785=>X"00",
7786=>X"00",
7787=>X"00",
7788=>X"00",
7789=>X"00",
7790=>X"00",
7791=>X"00",
7792=>X"00",
7793=>X"00",
7794=>X"00",
7795=>X"00",
7796=>X"00",
7797=>X"00",
7798=>X"00",
7799=>X"00",
7800=>X"00",
7801=>X"00",
7802=>X"00",
7803=>X"00",
7804=>X"00",
7805=>X"00",
7806=>X"00",
7807=>X"00",
7808=>X"00",
7809=>X"00",
7810=>X"00",
7811=>X"00",
7812=>X"00",
7813=>X"00",
7814=>X"00",
7815=>X"00",
7816=>X"00",
7817=>X"00",
7818=>X"00",
7819=>X"00",
7820=>X"00",
7821=>X"00",
7822=>X"00",
7823=>X"00",
7824=>X"00",
7825=>X"00",
7826=>X"00",
7827=>X"00",
7828=>X"00",
7829=>X"00",
7830=>X"00",
7831=>X"00",
7832=>X"00",
7833=>X"00",
7834=>X"00",
7835=>X"00",
7836=>X"00",
7837=>X"00",
7838=>X"00",
7839=>X"00",
7840=>X"00",
7841=>X"00",
7842=>X"00",
7843=>X"00",
7844=>X"00",
7845=>X"00",
7846=>X"00",
7847=>X"00",
7848=>X"00",
7849=>X"00",
7850=>X"00",
7851=>X"00",
7852=>X"00",
7853=>X"00",
7854=>X"00",
7855=>X"00",
7856=>X"00",
7857=>X"00",
7858=>X"00",
7859=>X"00",
7860=>X"00",
7861=>X"00",
7862=>X"00",
7863=>X"00",
7864=>X"00",
7865=>X"00",
7866=>X"00",
7867=>X"00",
7868=>X"00",
7869=>X"00",
7870=>X"00",
7871=>X"00",
7872=>X"00",
7873=>X"00",
7874=>X"00",
7875=>X"00",
7876=>X"00",
7877=>X"00",
7878=>X"00",
7879=>X"00",
7880=>X"00",
7881=>X"00",
7882=>X"00",
7883=>X"00",
7884=>X"00",
7885=>X"00",
7886=>X"00",
7887=>X"00",
7888=>X"00",
7889=>X"00",
7890=>X"00",
7891=>X"00",
7892=>X"00",
7893=>X"00",
7894=>X"00",
7895=>X"00",
7896=>X"00",
7897=>X"00",
7898=>X"00",
7899=>X"00",
7900=>X"00",
7901=>X"00",
7902=>X"00",
7903=>X"00",
7904=>X"00",
7905=>X"00",
7906=>X"00",
7907=>X"00",
7908=>X"00",
7909=>X"00",
7910=>X"00",
7911=>X"00",
7912=>X"00",
7913=>X"00",
7914=>X"00",
7915=>X"00",
7916=>X"00",
7917=>X"00",
7918=>X"00",
7919=>X"00",
7920=>X"00",
7921=>X"00",
7922=>X"00",
7923=>X"00",
7924=>X"00",
7925=>X"00",
7926=>X"00",
7927=>X"00",
7928=>X"00",
7929=>X"00",
7930=>X"00",
7931=>X"00",
7932=>X"00",
7933=>X"00",
7934=>X"00",
7935=>X"00",
7936=>X"15",
7937=>X"15",
7938=>X"15",
7939=>X"15",
7940=>X"15",
7941=>X"15",
7942=>X"15",
7943=>X"15",
7944=>X"14",
7945=>X"14",
7946=>X"14",
7947=>X"14",
7948=>X"14",
7949=>X"14",
7950=>X"14",
7951=>X"14",
7952=>X"14",
7953=>X"14",
7954=>X"14",
7955=>X"14",
7956=>X"14",
7957=>X"14",
7958=>X"15",
7959=>X"15",
7960=>X"15",
7961=>X"15",
7962=>X"15",
7963=>X"15",
7964=>X"15",
7965=>X"15",
7966=>X"15",
7967=>X"15",
7968=>X"15",
7969=>X"15",
7970=>X"19",
7971=>X"29",
7972=>X"29",
7973=>X"29",
7974=>X"19",
7975=>X"19",
7976=>X"19",
7977=>X"19",
7978=>X"19",
7979=>X"19",
7980=>X"19",
7981=>X"19",
7982=>X"19",
7983=>X"19",
7984=>X"19",
7985=>X"19",
7986=>X"19",
7987=>X"19",
7988=>X"19",
7989=>X"2A",
7990=>X"1A",
7991=>X"1A",
7992=>X"2A",
7993=>X"1A",
7994=>X"1A",
7995=>X"1A",
7996=>X"26",
7997=>X"26",
7998=>X"27",
7999=>X"27",
8000=>X"26",
8001=>X"15",
8002=>X"15",
8003=>X"15",
8004=>X"15",
8005=>X"15",
8006=>X"15",
8007=>X"15",
8008=>X"15",
8009=>X"15",
8010=>X"15",
8011=>X"15",
8012=>X"15",
8013=>X"15",
8014=>X"15",
8015=>X"15",
8016=>X"15",
8017=>X"15",
8018=>X"15",
8019=>X"15",
8020=>X"15",
8021=>X"15",
8022=>X"15",
8023=>X"15",
8024=>X"15",
8025=>X"15",
8026=>X"15",
8027=>X"15",
8028=>X"15",
8029=>X"15",
8030=>X"15",
8031=>X"15",
8032=>X"15",
8033=>X"15",
8034=>X"15",
8035=>X"15",
8036=>X"00",
8037=>X"00",
8038=>X"00",
8039=>X"00",
8040=>X"00",
8041=>X"00",
8042=>X"00",
8043=>X"00",
8044=>X"00",
8045=>X"00",
8046=>X"00",
8047=>X"00",
8048=>X"00",
8049=>X"00",
8050=>X"00",
8051=>X"00",
8052=>X"00",
8053=>X"00",
8054=>X"00",
8055=>X"00",
8056=>X"00",
8057=>X"00",
8058=>X"00",
8059=>X"00",
8060=>X"00",
8061=>X"00",
8062=>X"00",
8063=>X"00",
8064=>X"00",
8065=>X"00",
8066=>X"00",
8067=>X"00",
8068=>X"00",
8069=>X"00",
8070=>X"00",
8071=>X"00",
8072=>X"00",
8073=>X"00",
8074=>X"00",
8075=>X"00",
8076=>X"00",
8077=>X"00",
8078=>X"00",
8079=>X"00",
8080=>X"00",
8081=>X"00",
8082=>X"00",
8083=>X"00",
8084=>X"00",
8085=>X"00",
8086=>X"00",
8087=>X"00",
8088=>X"00",
8089=>X"00",
8090=>X"00",
8091=>X"00",
8092=>X"00",
8093=>X"00",
8094=>X"00",
8095=>X"00",
8096=>X"00",
8097=>X"00",
8098=>X"00",
8099=>X"00",
8100=>X"00",
8101=>X"00",
8102=>X"00",
8103=>X"00",
8104=>X"00",
8105=>X"00",
8106=>X"00",
8107=>X"00",
8108=>X"00",
8109=>X"00",
8110=>X"00",
8111=>X"00",
8112=>X"00",
8113=>X"00",
8114=>X"00",
8115=>X"00",
8116=>X"00",
8117=>X"00",
8118=>X"00",
8119=>X"00",
8120=>X"00",
8121=>X"00",
8122=>X"00",
8123=>X"00",
8124=>X"00",
8125=>X"00",
8126=>X"00",
8127=>X"00",
8128=>X"00",
8129=>X"00",
8130=>X"00",
8131=>X"00",
8132=>X"00",
8133=>X"00",
8134=>X"00",
8135=>X"00",
8136=>X"00",
8137=>X"00",
8138=>X"00",
8139=>X"00",
8140=>X"00",
8141=>X"00",
8142=>X"00",
8143=>X"00",
8144=>X"00",
8145=>X"00",
8146=>X"00",
8147=>X"00",
8148=>X"00",
8149=>X"00",
8150=>X"00",
8151=>X"00",
8152=>X"00",
8153=>X"00",
8154=>X"00",
8155=>X"00",
8156=>X"00",
8157=>X"00",
8158=>X"00",
8159=>X"00",
8160=>X"00",
8161=>X"00",
8162=>X"00",
8163=>X"00",
8164=>X"00",
8165=>X"00",
8166=>X"00",
8167=>X"00",
8168=>X"00",
8169=>X"00",
8170=>X"00",
8171=>X"00",
8172=>X"00",
8173=>X"00",
8174=>X"00",
8175=>X"00",
8176=>X"00",
8177=>X"00",
8178=>X"00",
8179=>X"00",
8180=>X"00",
8181=>X"00",
8182=>X"00",
8183=>X"00",
8184=>X"00",
8185=>X"00",
8186=>X"00",
8187=>X"00",
8188=>X"00",
8189=>X"00",
8190=>X"00",
8191=>X"00",
8192=>X"15",
8193=>X"15",
8194=>X"15",
8195=>X"15",
8196=>X"15",
8197=>X"15",
8198=>X"15",
8199=>X"15",
8200=>X"15",
8201=>X"15",
8202=>X"14",
8203=>X"14",
8204=>X"14",
8205=>X"14",
8206=>X"14",
8207=>X"14",
8208=>X"14",
8209=>X"14",
8210=>X"14",
8211=>X"14",
8212=>X"14",
8213=>X"14",
8214=>X"15",
8215=>X"15",
8216=>X"15",
8217=>X"15",
8218=>X"15",
8219=>X"15",
8220=>X"15",
8221=>X"15",
8222=>X"15",
8223=>X"15",
8224=>X"15",
8225=>X"15",
8226=>X"29",
8227=>X"29",
8228=>X"29",
8229=>X"19",
8230=>X"19",
8231=>X"19",
8232=>X"19",
8233=>X"19",
8234=>X"19",
8235=>X"19",
8236=>X"19",
8237=>X"19",
8238=>X"19",
8239=>X"19",
8240=>X"19",
8241=>X"19",
8242=>X"19",
8243=>X"19",
8244=>X"1A",
8245=>X"1A",
8246=>X"1A",
8247=>X"19",
8248=>X"1A",
8249=>X"1A",
8250=>X"1A",
8251=>X"19",
8252=>X"15",
8253=>X"16",
8254=>X"27",
8255=>X"27",
8256=>X"27",
8257=>X"26",
8258=>X"15",
8259=>X"15",
8260=>X"15",
8261=>X"15",
8262=>X"15",
8263=>X"15",
8264=>X"15",
8265=>X"15",
8266=>X"15",
8267=>X"15",
8268=>X"15",
8269=>X"15",
8270=>X"15",
8271=>X"15",
8272=>X"15",
8273=>X"15",
8274=>X"15",
8275=>X"15",
8276=>X"15",
8277=>X"15",
8278=>X"15",
8279=>X"15",
8280=>X"15",
8281=>X"15",
8282=>X"15",
8283=>X"15",
8284=>X"15",
8285=>X"15",
8286=>X"15",
8287=>X"15",
8288=>X"19",
8289=>X"19",
8290=>X"19",
8291=>X"19",
8292=>X"00",
8293=>X"00",
8294=>X"00",
8295=>X"00",
8296=>X"00",
8297=>X"00",
8298=>X"00",
8299=>X"00",
8300=>X"00",
8301=>X"00",
8302=>X"00",
8303=>X"00",
8304=>X"00",
8305=>X"00",
8306=>X"00",
8307=>X"00",
8308=>X"00",
8309=>X"00",
8310=>X"00",
8311=>X"00",
8312=>X"00",
8313=>X"00",
8314=>X"00",
8315=>X"00",
8316=>X"00",
8317=>X"00",
8318=>X"00",
8319=>X"00",
8320=>X"00",
8321=>X"00",
8322=>X"00",
8323=>X"00",
8324=>X"00",
8325=>X"00",
8326=>X"00",
8327=>X"00",
8328=>X"00",
8329=>X"00",
8330=>X"00",
8331=>X"00",
8332=>X"00",
8333=>X"00",
8334=>X"00",
8335=>X"00",
8336=>X"00",
8337=>X"00",
8338=>X"00",
8339=>X"00",
8340=>X"00",
8341=>X"00",
8342=>X"00",
8343=>X"00",
8344=>X"00",
8345=>X"00",
8346=>X"00",
8347=>X"00",
8348=>X"00",
8349=>X"00",
8350=>X"00",
8351=>X"00",
8352=>X"00",
8353=>X"00",
8354=>X"00",
8355=>X"00",
8356=>X"00",
8357=>X"00",
8358=>X"00",
8359=>X"00",
8360=>X"00",
8361=>X"00",
8362=>X"00",
8363=>X"00",
8364=>X"00",
8365=>X"00",
8366=>X"00",
8367=>X"00",
8368=>X"00",
8369=>X"00",
8370=>X"00",
8371=>X"00",
8372=>X"00",
8373=>X"00",
8374=>X"00",
8375=>X"00",
8376=>X"00",
8377=>X"00",
8378=>X"00",
8379=>X"00",
8380=>X"00",
8381=>X"00",
8382=>X"00",
8383=>X"00",
8384=>X"00",
8385=>X"00",
8386=>X"00",
8387=>X"00",
8388=>X"00",
8389=>X"00",
8390=>X"00",
8391=>X"00",
8392=>X"00",
8393=>X"00",
8394=>X"00",
8395=>X"00",
8396=>X"00",
8397=>X"00",
8398=>X"00",
8399=>X"00",
8400=>X"00",
8401=>X"00",
8402=>X"00",
8403=>X"00",
8404=>X"00",
8405=>X"00",
8406=>X"00",
8407=>X"00",
8408=>X"00",
8409=>X"00",
8410=>X"00",
8411=>X"00",
8412=>X"00",
8413=>X"00",
8414=>X"00",
8415=>X"00",
8416=>X"00",
8417=>X"00",
8418=>X"00",
8419=>X"00",
8420=>X"00",
8421=>X"00",
8422=>X"00",
8423=>X"00",
8424=>X"00",
8425=>X"00",
8426=>X"00",
8427=>X"00",
8428=>X"00",
8429=>X"00",
8430=>X"00",
8431=>X"00",
8432=>X"00",
8433=>X"00",
8434=>X"00",
8435=>X"00",
8436=>X"00",
8437=>X"00",
8438=>X"00",
8439=>X"00",
8440=>X"00",
8441=>X"00",
8442=>X"00",
8443=>X"00",
8444=>X"00",
8445=>X"00",
8446=>X"00",
8447=>X"00",
8448=>X"15",
8449=>X"15",
8450=>X"15",
8451=>X"15",
8452=>X"15",
8453=>X"15",
8454=>X"15",
8455=>X"15",
8456=>X"15",
8457=>X"15",
8458=>X"14",
8459=>X"15",
8460=>X"15",
8461=>X"15",
8462=>X"15",
8463=>X"15",
8464=>X"15",
8465=>X"15",
8466=>X"14",
8467=>X"14",
8468=>X"14",
8469=>X"14",
8470=>X"15",
8471=>X"15",
8472=>X"15",
8473=>X"15",
8474=>X"15",
8475=>X"15",
8476=>X"15",
8477=>X"15",
8478=>X"15",
8479=>X"15",
8480=>X"15",
8481=>X"29",
8482=>X"29",
8483=>X"29",
8484=>X"29",
8485=>X"19",
8486=>X"19",
8487=>X"19",
8488=>X"19",
8489=>X"19",
8490=>X"19",
8491=>X"19",
8492=>X"19",
8493=>X"19",
8494=>X"19",
8495=>X"19",
8496=>X"19",
8497=>X"19",
8498=>X"19",
8499=>X"19",
8500=>X"19",
8501=>X"1A",
8502=>X"19",
8503=>X"19",
8504=>X"19",
8505=>X"1A",
8506=>X"2A",
8507=>X"19",
8508=>X"15",
8509=>X"15",
8510=>X"16",
8511=>X"27",
8512=>X"27",
8513=>X"26",
8514=>X"15",
8515=>X"15",
8516=>X"15",
8517=>X"15",
8518=>X"15",
8519=>X"15",
8520=>X"15",
8521=>X"15",
8522=>X"15",
8523=>X"15",
8524=>X"15",
8525=>X"15",
8526=>X"15",
8527=>X"15",
8528=>X"15",
8529=>X"15",
8530=>X"15",
8531=>X"15",
8532=>X"15",
8533=>X"15",
8534=>X"15",
8535=>X"15",
8536=>X"15",
8537=>X"15",
8538=>X"15",
8539=>X"15",
8540=>X"15",
8541=>X"15",
8542=>X"15",
8543=>X"15",
8544=>X"19",
8545=>X"15",
8546=>X"19",
8547=>X"15",
8548=>X"00",
8549=>X"00",
8550=>X"00",
8551=>X"00",
8552=>X"00",
8553=>X"00",
8554=>X"00",
8555=>X"00",
8556=>X"00",
8557=>X"00",
8558=>X"00",
8559=>X"00",
8560=>X"00",
8561=>X"00",
8562=>X"00",
8563=>X"00",
8564=>X"00",
8565=>X"00",
8566=>X"00",
8567=>X"00",
8568=>X"00",
8569=>X"00",
8570=>X"00",
8571=>X"00",
8572=>X"00",
8573=>X"00",
8574=>X"00",
8575=>X"00",
8576=>X"00",
8577=>X"00",
8578=>X"00",
8579=>X"00",
8580=>X"00",
8581=>X"00",
8582=>X"00",
8583=>X"00",
8584=>X"00",
8585=>X"00",
8586=>X"00",
8587=>X"00",
8588=>X"00",
8589=>X"00",
8590=>X"00",
8591=>X"00",
8592=>X"00",
8593=>X"00",
8594=>X"00",
8595=>X"00",
8596=>X"00",
8597=>X"00",
8598=>X"00",
8599=>X"00",
8600=>X"00",
8601=>X"00",
8602=>X"00",
8603=>X"00",
8604=>X"00",
8605=>X"00",
8606=>X"00",
8607=>X"00",
8608=>X"00",
8609=>X"00",
8610=>X"00",
8611=>X"00",
8612=>X"00",
8613=>X"00",
8614=>X"00",
8615=>X"00",
8616=>X"00",
8617=>X"00",
8618=>X"00",
8619=>X"00",
8620=>X"00",
8621=>X"00",
8622=>X"00",
8623=>X"00",
8624=>X"00",
8625=>X"00",
8626=>X"00",
8627=>X"00",
8628=>X"00",
8629=>X"00",
8630=>X"00",
8631=>X"00",
8632=>X"00",
8633=>X"00",
8634=>X"00",
8635=>X"00",
8636=>X"00",
8637=>X"00",
8638=>X"00",
8639=>X"00",
8640=>X"00",
8641=>X"00",
8642=>X"00",
8643=>X"00",
8644=>X"00",
8645=>X"00",
8646=>X"00",
8647=>X"00",
8648=>X"00",
8649=>X"00",
8650=>X"00",
8651=>X"00",
8652=>X"00",
8653=>X"00",
8654=>X"00",
8655=>X"00",
8656=>X"00",
8657=>X"00",
8658=>X"00",
8659=>X"00",
8660=>X"00",
8661=>X"00",
8662=>X"00",
8663=>X"00",
8664=>X"00",
8665=>X"00",
8666=>X"00",
8667=>X"00",
8668=>X"00",
8669=>X"00",
8670=>X"00",
8671=>X"00",
8672=>X"00",
8673=>X"00",
8674=>X"00",
8675=>X"00",
8676=>X"00",
8677=>X"00",
8678=>X"00",
8679=>X"00",
8680=>X"00",
8681=>X"00",
8682=>X"00",
8683=>X"00",
8684=>X"00",
8685=>X"00",
8686=>X"00",
8687=>X"00",
8688=>X"00",
8689=>X"00",
8690=>X"00",
8691=>X"00",
8692=>X"00",
8693=>X"00",
8694=>X"00",
8695=>X"00",
8696=>X"00",
8697=>X"00",
8698=>X"00",
8699=>X"00",
8700=>X"00",
8701=>X"00",
8702=>X"00",
8703=>X"00",
8704=>X"15",
8705=>X"15",
8706=>X"15",
8707=>X"15",
8708=>X"15",
8709=>X"15",
8710=>X"15",
8711=>X"15",
8712=>X"15",
8713=>X"15",
8714=>X"14",
8715=>X"15",
8716=>X"15",
8717=>X"15",
8718=>X"15",
8719=>X"15",
8720=>X"15",
8721=>X"15",
8722=>X"15",
8723=>X"15",
8724=>X"14",
8725=>X"14",
8726=>X"15",
8727=>X"15",
8728=>X"15",
8729=>X"15",
8730=>X"15",
8731=>X"15",
8732=>X"15",
8733=>X"15",
8734=>X"15",
8735=>X"15",
8736=>X"29",
8737=>X"29",
8738=>X"29",
8739=>X"19",
8740=>X"19",
8741=>X"19",
8742=>X"29",
8743=>X"19",
8744=>X"19",
8745=>X"19",
8746=>X"19",
8747=>X"19",
8748=>X"19",
8749=>X"19",
8750=>X"19",
8751=>X"19",
8752=>X"19",
8753=>X"19",
8754=>X"19",
8755=>X"19",
8756=>X"19",
8757=>X"19",
8758=>X"19",
8759=>X"19",
8760=>X"19",
8761=>X"2A",
8762=>X"2E",
8763=>X"2A",
8764=>X"15",
8765=>X"15",
8766=>X"16",
8767=>X"26",
8768=>X"26",
8769=>X"26",
8770=>X"15",
8771=>X"15",
8772=>X"15",
8773=>X"15",
8774=>X"15",
8775=>X"15",
8776=>X"15",
8777=>X"15",
8778=>X"15",
8779=>X"15",
8780=>X"15",
8781=>X"15",
8782=>X"15",
8783=>X"15",
8784=>X"15",
8785=>X"15",
8786=>X"15",
8787=>X"15",
8788=>X"15",
8789=>X"15",
8790=>X"15",
8791=>X"15",
8792=>X"15",
8793=>X"15",
8794=>X"15",
8795=>X"15",
8796=>X"15",
8797=>X"19",
8798=>X"15",
8799=>X"15",
8800=>X"15",
8801=>X"15",
8802=>X"15",
8803=>X"15",
8804=>X"00",
8805=>X"00",
8806=>X"00",
8807=>X"00",
8808=>X"00",
8809=>X"00",
8810=>X"00",
8811=>X"00",
8812=>X"00",
8813=>X"00",
8814=>X"00",
8815=>X"00",
8816=>X"00",
8817=>X"00",
8818=>X"00",
8819=>X"00",
8820=>X"00",
8821=>X"00",
8822=>X"00",
8823=>X"00",
8824=>X"00",
8825=>X"00",
8826=>X"00",
8827=>X"00",
8828=>X"00",
8829=>X"00",
8830=>X"00",
8831=>X"00",
8832=>X"00",
8833=>X"00",
8834=>X"00",
8835=>X"00",
8836=>X"00",
8837=>X"00",
8838=>X"00",
8839=>X"00",
8840=>X"00",
8841=>X"00",
8842=>X"00",
8843=>X"00",
8844=>X"00",
8845=>X"00",
8846=>X"00",
8847=>X"00",
8848=>X"00",
8849=>X"00",
8850=>X"00",
8851=>X"00",
8852=>X"00",
8853=>X"00",
8854=>X"00",
8855=>X"00",
8856=>X"00",
8857=>X"00",
8858=>X"00",
8859=>X"00",
8860=>X"00",
8861=>X"00",
8862=>X"00",
8863=>X"00",
8864=>X"00",
8865=>X"00",
8866=>X"00",
8867=>X"00",
8868=>X"00",
8869=>X"00",
8870=>X"00",
8871=>X"00",
8872=>X"00",
8873=>X"00",
8874=>X"00",
8875=>X"00",
8876=>X"00",
8877=>X"00",
8878=>X"00",
8879=>X"00",
8880=>X"00",
8881=>X"00",
8882=>X"00",
8883=>X"00",
8884=>X"00",
8885=>X"00",
8886=>X"00",
8887=>X"00",
8888=>X"00",
8889=>X"00",
8890=>X"00",
8891=>X"00",
8892=>X"00",
8893=>X"00",
8894=>X"00",
8895=>X"00",
8896=>X"00",
8897=>X"00",
8898=>X"00",
8899=>X"00",
8900=>X"00",
8901=>X"00",
8902=>X"00",
8903=>X"00",
8904=>X"00",
8905=>X"00",
8906=>X"00",
8907=>X"00",
8908=>X"00",
8909=>X"00",
8910=>X"00",
8911=>X"00",
8912=>X"00",
8913=>X"00",
8914=>X"00",
8915=>X"00",
8916=>X"00",
8917=>X"00",
8918=>X"00",
8919=>X"00",
8920=>X"00",
8921=>X"00",
8922=>X"00",
8923=>X"00",
8924=>X"00",
8925=>X"00",
8926=>X"00",
8927=>X"00",
8928=>X"00",
8929=>X"00",
8930=>X"00",
8931=>X"00",
8932=>X"00",
8933=>X"00",
8934=>X"00",
8935=>X"00",
8936=>X"00",
8937=>X"00",
8938=>X"00",
8939=>X"00",
8940=>X"00",
8941=>X"00",
8942=>X"00",
8943=>X"00",
8944=>X"00",
8945=>X"00",
8946=>X"00",
8947=>X"00",
8948=>X"00",
8949=>X"00",
8950=>X"00",
8951=>X"00",
8952=>X"00",
8953=>X"00",
8954=>X"00",
8955=>X"00",
8956=>X"00",
8957=>X"00",
8958=>X"00",
8959=>X"00",
8960=>X"15",
8961=>X"15",
8962=>X"15",
8963=>X"15",
8964=>X"15",
8965=>X"15",
8966=>X"15",
8967=>X"15",
8968=>X"15",
8969=>X"15",
8970=>X"15",
8971=>X"15",
8972=>X"15",
8973=>X"15",
8974=>X"15",
8975=>X"15",
8976=>X"15",
8977=>X"15",
8978=>X"15",
8979=>X"15",
8980=>X"15",
8981=>X"15",
8982=>X"15",
8983=>X"15",
8984=>X"15",
8985=>X"15",
8986=>X"15",
8987=>X"15",
8988=>X"15",
8989=>X"15",
8990=>X"15",
8991=>X"19",
8992=>X"29",
8993=>X"29",
8994=>X"29",
8995=>X"29",
8996=>X"19",
8997=>X"19",
8998=>X"29",
8999=>X"19",
9000=>X"19",
9001=>X"19",
9002=>X"19",
9003=>X"19",
9004=>X"19",
9005=>X"19",
9006=>X"19",
9007=>X"19",
9008=>X"19",
9009=>X"19",
9010=>X"19",
9011=>X"19",
9012=>X"19",
9013=>X"19",
9014=>X"29",
9015=>X"2A",
9016=>X"2A",
9017=>X"3E",
9018=>X"3F",
9019=>X"2B",
9020=>X"2A",
9021=>X"25",
9022=>X"26",
9023=>X"27",
9024=>X"16",
9025=>X"26",
9026=>X"16",
9027=>X"15",
9028=>X"15",
9029=>X"15",
9030=>X"15",
9031=>X"15",
9032=>X"15",
9033=>X"15",
9034=>X"15",
9035=>X"15",
9036=>X"15",
9037=>X"15",
9038=>X"15",
9039=>X"15",
9040=>X"15",
9041=>X"15",
9042=>X"15",
9043=>X"15",
9044=>X"19",
9045=>X"15",
9046=>X"19",
9047=>X"15",
9048=>X"15",
9049=>X"15",
9050=>X"15",
9051=>X"15",
9052=>X"15",
9053=>X"19",
9054=>X"15",
9055=>X"15",
9056=>X"15",
9057=>X"15",
9058=>X"15",
9059=>X"15",
9060=>X"00",
9061=>X"00",
9062=>X"00",
9063=>X"00",
9064=>X"00",
9065=>X"00",
9066=>X"00",
9067=>X"00",
9068=>X"00",
9069=>X"00",
9070=>X"00",
9071=>X"00",
9072=>X"00",
9073=>X"00",
9074=>X"00",
9075=>X"00",
9076=>X"00",
9077=>X"00",
9078=>X"00",
9079=>X"00",
9080=>X"00",
9081=>X"00",
9082=>X"00",
9083=>X"00",
9084=>X"00",
9085=>X"00",
9086=>X"00",
9087=>X"00",
9088=>X"00",
9089=>X"00",
9090=>X"00",
9091=>X"00",
9092=>X"00",
9093=>X"00",
9094=>X"00",
9095=>X"00",
9096=>X"00",
9097=>X"00",
9098=>X"00",
9099=>X"00",
9100=>X"00",
9101=>X"00",
9102=>X"00",
9103=>X"00",
9104=>X"00",
9105=>X"00",
9106=>X"00",
9107=>X"00",
9108=>X"00",
9109=>X"00",
9110=>X"00",
9111=>X"00",
9112=>X"00",
9113=>X"00",
9114=>X"00",
9115=>X"00",
9116=>X"00",
9117=>X"00",
9118=>X"00",
9119=>X"00",
9120=>X"00",
9121=>X"00",
9122=>X"00",
9123=>X"00",
9124=>X"00",
9125=>X"00",
9126=>X"00",
9127=>X"00",
9128=>X"00",
9129=>X"00",
9130=>X"00",
9131=>X"00",
9132=>X"00",
9133=>X"00",
9134=>X"00",
9135=>X"00",
9136=>X"00",
9137=>X"00",
9138=>X"00",
9139=>X"00",
9140=>X"00",
9141=>X"00",
9142=>X"00",
9143=>X"00",
9144=>X"00",
9145=>X"00",
9146=>X"00",
9147=>X"00",
9148=>X"00",
9149=>X"00",
9150=>X"00",
9151=>X"00",
9152=>X"00",
9153=>X"00",
9154=>X"00",
9155=>X"00",
9156=>X"00",
9157=>X"00",
9158=>X"00",
9159=>X"00",
9160=>X"00",
9161=>X"00",
9162=>X"00",
9163=>X"00",
9164=>X"00",
9165=>X"00",
9166=>X"00",
9167=>X"00",
9168=>X"00",
9169=>X"00",
9170=>X"00",
9171=>X"00",
9172=>X"00",
9173=>X"00",
9174=>X"00",
9175=>X"00",
9176=>X"00",
9177=>X"00",
9178=>X"00",
9179=>X"00",
9180=>X"00",
9181=>X"00",
9182=>X"00",
9183=>X"00",
9184=>X"00",
9185=>X"00",
9186=>X"00",
9187=>X"00",
9188=>X"00",
9189=>X"00",
9190=>X"00",
9191=>X"00",
9192=>X"00",
9193=>X"00",
9194=>X"00",
9195=>X"00",
9196=>X"00",
9197=>X"00",
9198=>X"00",
9199=>X"00",
9200=>X"00",
9201=>X"00",
9202=>X"00",
9203=>X"00",
9204=>X"00",
9205=>X"00",
9206=>X"00",
9207=>X"00",
9208=>X"00",
9209=>X"00",
9210=>X"00",
9211=>X"00",
9212=>X"00",
9213=>X"00",
9214=>X"00",
9215=>X"00",
9216=>X"15",
9217=>X"15",
9218=>X"15",
9219=>X"15",
9220=>X"15",
9221=>X"15",
9222=>X"15",
9223=>X"15",
9224=>X"15",
9225=>X"15",
9226=>X"15",
9227=>X"15",
9228=>X"15",
9229=>X"15",
9230=>X"15",
9231=>X"15",
9232=>X"15",
9233=>X"15",
9234=>X"15",
9235=>X"15",
9236=>X"15",
9237=>X"15",
9238=>X"15",
9239=>X"15",
9240=>X"15",
9241=>X"15",
9242=>X"15",
9243=>X"15",
9244=>X"15",
9245=>X"15",
9246=>X"29",
9247=>X"2D",
9248=>X"2D",
9249=>X"29",
9250=>X"29",
9251=>X"29",
9252=>X"19",
9253=>X"19",
9254=>X"19",
9255=>X"19",
9256=>X"19",
9257=>X"19",
9258=>X"19",
9259=>X"19",
9260=>X"19",
9261=>X"19",
9262=>X"19",
9263=>X"19",
9264=>X"19",
9265=>X"19",
9266=>X"19",
9267=>X"19",
9268=>X"19",
9269=>X"2A",
9270=>X"3E",
9271=>X"3E",
9272=>X"3E",
9273=>X"3E",
9274=>X"3F",
9275=>X"3A",
9276=>X"2A",
9277=>X"29",
9278=>X"26",
9279=>X"17",
9280=>X"16",
9281=>X"16",
9282=>X"26",
9283=>X"16",
9284=>X"15",
9285=>X"15",
9286=>X"15",
9287=>X"15",
9288=>X"15",
9289=>X"15",
9290=>X"15",
9291=>X"15",
9292=>X"15",
9293=>X"15",
9294=>X"15",
9295=>X"15",
9296=>X"15",
9297=>X"19",
9298=>X"15",
9299=>X"15",
9300=>X"19",
9301=>X"15",
9302=>X"19",
9303=>X"15",
9304=>X"15",
9305=>X"15",
9306=>X"15",
9307=>X"15",
9308=>X"15",
9309=>X"15",
9310=>X"15",
9311=>X"15",
9312=>X"15",
9313=>X"15",
9314=>X"15",
9315=>X"15",
9316=>X"00",
9317=>X"00",
9318=>X"00",
9319=>X"00",
9320=>X"00",
9321=>X"00",
9322=>X"00",
9323=>X"00",
9324=>X"00",
9325=>X"00",
9326=>X"00",
9327=>X"00",
9328=>X"00",
9329=>X"00",
9330=>X"00",
9331=>X"00",
9332=>X"00",
9333=>X"00",
9334=>X"00",
9335=>X"00",
9336=>X"00",
9337=>X"00",
9338=>X"00",
9339=>X"00",
9340=>X"00",
9341=>X"00",
9342=>X"00",
9343=>X"00",
9344=>X"00",
9345=>X"00",
9346=>X"00",
9347=>X"00",
9348=>X"00",
9349=>X"00",
9350=>X"00",
9351=>X"00",
9352=>X"00",
9353=>X"00",
9354=>X"00",
9355=>X"00",
9356=>X"00",
9357=>X"00",
9358=>X"00",
9359=>X"00",
9360=>X"00",
9361=>X"00",
9362=>X"00",
9363=>X"00",
9364=>X"00",
9365=>X"00",
9366=>X"00",
9367=>X"00",
9368=>X"00",
9369=>X"00",
9370=>X"00",
9371=>X"00",
9372=>X"00",
9373=>X"00",
9374=>X"00",
9375=>X"00",
9376=>X"00",
9377=>X"00",
9378=>X"00",
9379=>X"00",
9380=>X"00",
9381=>X"00",
9382=>X"00",
9383=>X"00",
9384=>X"00",
9385=>X"00",
9386=>X"00",
9387=>X"00",
9388=>X"00",
9389=>X"00",
9390=>X"00",
9391=>X"00",
9392=>X"00",
9393=>X"00",
9394=>X"00",
9395=>X"00",
9396=>X"00",
9397=>X"00",
9398=>X"00",
9399=>X"00",
9400=>X"00",
9401=>X"00",
9402=>X"00",
9403=>X"00",
9404=>X"00",
9405=>X"00",
9406=>X"00",
9407=>X"00",
9408=>X"00",
9409=>X"00",
9410=>X"00",
9411=>X"00",
9412=>X"00",
9413=>X"00",
9414=>X"00",
9415=>X"00",
9416=>X"00",
9417=>X"00",
9418=>X"00",
9419=>X"00",
9420=>X"00",
9421=>X"00",
9422=>X"00",
9423=>X"00",
9424=>X"00",
9425=>X"00",
9426=>X"00",
9427=>X"00",
9428=>X"00",
9429=>X"00",
9430=>X"00",
9431=>X"00",
9432=>X"00",
9433=>X"00",
9434=>X"00",
9435=>X"00",
9436=>X"00",
9437=>X"00",
9438=>X"00",
9439=>X"00",
9440=>X"00",
9441=>X"00",
9442=>X"00",
9443=>X"00",
9444=>X"00",
9445=>X"00",
9446=>X"00",
9447=>X"00",
9448=>X"00",
9449=>X"00",
9450=>X"00",
9451=>X"00",
9452=>X"00",
9453=>X"00",
9454=>X"00",
9455=>X"00",
9456=>X"00",
9457=>X"00",
9458=>X"00",
9459=>X"00",
9460=>X"00",
9461=>X"00",
9462=>X"00",
9463=>X"00",
9464=>X"00",
9465=>X"00",
9466=>X"00",
9467=>X"00",
9468=>X"00",
9469=>X"00",
9470=>X"00",
9471=>X"00",
9472=>X"15",
9473=>X"15",
9474=>X"15",
9475=>X"15",
9476=>X"15",
9477=>X"15",
9478=>X"15",
9479=>X"15",
9480=>X"15",
9481=>X"15",
9482=>X"15",
9483=>X"15",
9484=>X"15",
9485=>X"15",
9486=>X"15",
9487=>X"15",
9488=>X"15",
9489=>X"15",
9490=>X"15",
9491=>X"15",
9492=>X"15",
9493=>X"15",
9494=>X"15",
9495=>X"15",
9496=>X"15",
9497=>X"15",
9498=>X"15",
9499=>X"15",
9500=>X"15",
9501=>X"15",
9502=>X"2E",
9503=>X"2E",
9504=>X"2E",
9505=>X"29",
9506=>X"1A",
9507=>X"29",
9508=>X"19",
9509=>X"19",
9510=>X"19",
9511=>X"19",
9512=>X"19",
9513=>X"19",
9514=>X"19",
9515=>X"19",
9516=>X"19",
9517=>X"19",
9518=>X"19",
9519=>X"19",
9520=>X"19",
9521=>X"19",
9522=>X"2A",
9523=>X"2A",
9524=>X"2A",
9525=>X"2A",
9526=>X"3E",
9527=>X"3E",
9528=>X"3E",
9529=>X"3E",
9530=>X"3A",
9531=>X"2A",
9532=>X"2A",
9533=>X"29",
9534=>X"26",
9535=>X"26",
9536=>X"16",
9537=>X"16",
9538=>X"26",
9539=>X"16",
9540=>X"15",
9541=>X"15",
9542=>X"15",
9543=>X"15",
9544=>X"15",
9545=>X"15",
9546=>X"15",
9547=>X"15",
9548=>X"15",
9549=>X"15",
9550=>X"15",
9551=>X"19",
9552=>X"15",
9553=>X"19",
9554=>X"15",
9555=>X"15",
9556=>X"15",
9557=>X"15",
9558=>X"15",
9559=>X"15",
9560=>X"15",
9561=>X"15",
9562=>X"15",
9563=>X"15",
9564=>X"15",
9565=>X"15",
9566=>X"15",
9567=>X"15",
9568=>X"15",
9569=>X"15",
9570=>X"15",
9571=>X"15",
9572=>X"00",
9573=>X"00",
9574=>X"00",
9575=>X"00",
9576=>X"00",
9577=>X"00",
9578=>X"00",
9579=>X"00",
9580=>X"00",
9581=>X"00",
9582=>X"00",
9583=>X"00",
9584=>X"00",
9585=>X"00",
9586=>X"00",
9587=>X"00",
9588=>X"00",
9589=>X"00",
9590=>X"00",
9591=>X"00",
9592=>X"00",
9593=>X"00",
9594=>X"00",
9595=>X"00",
9596=>X"00",
9597=>X"00",
9598=>X"00",
9599=>X"00",
9600=>X"00",
9601=>X"00",
9602=>X"00",
9603=>X"00",
9604=>X"00",
9605=>X"00",
9606=>X"00",
9607=>X"00",
9608=>X"00",
9609=>X"00",
9610=>X"00",
9611=>X"00",
9612=>X"00",
9613=>X"00",
9614=>X"00",
9615=>X"00",
9616=>X"00",
9617=>X"00",
9618=>X"00",
9619=>X"00",
9620=>X"00",
9621=>X"00",
9622=>X"00",
9623=>X"00",
9624=>X"00",
9625=>X"00",
9626=>X"00",
9627=>X"00",
9628=>X"00",
9629=>X"00",
9630=>X"00",
9631=>X"00",
9632=>X"00",
9633=>X"00",
9634=>X"00",
9635=>X"00",
9636=>X"00",
9637=>X"00",
9638=>X"00",
9639=>X"00",
9640=>X"00",
9641=>X"00",
9642=>X"00",
9643=>X"00",
9644=>X"00",
9645=>X"00",
9646=>X"00",
9647=>X"00",
9648=>X"00",
9649=>X"00",
9650=>X"00",
9651=>X"00",
9652=>X"00",
9653=>X"00",
9654=>X"00",
9655=>X"00",
9656=>X"00",
9657=>X"00",
9658=>X"00",
9659=>X"00",
9660=>X"00",
9661=>X"00",
9662=>X"00",
9663=>X"00",
9664=>X"00",
9665=>X"00",
9666=>X"00",
9667=>X"00",
9668=>X"00",
9669=>X"00",
9670=>X"00",
9671=>X"00",
9672=>X"00",
9673=>X"00",
9674=>X"00",
9675=>X"00",
9676=>X"00",
9677=>X"00",
9678=>X"00",
9679=>X"00",
9680=>X"00",
9681=>X"00",
9682=>X"00",
9683=>X"00",
9684=>X"00",
9685=>X"00",
9686=>X"00",
9687=>X"00",
9688=>X"00",
9689=>X"00",
9690=>X"00",
9691=>X"00",
9692=>X"00",
9693=>X"00",
9694=>X"00",
9695=>X"00",
9696=>X"00",
9697=>X"00",
9698=>X"00",
9699=>X"00",
9700=>X"00",
9701=>X"00",
9702=>X"00",
9703=>X"00",
9704=>X"00",
9705=>X"00",
9706=>X"00",
9707=>X"00",
9708=>X"00",
9709=>X"00",
9710=>X"00",
9711=>X"00",
9712=>X"00",
9713=>X"00",
9714=>X"00",
9715=>X"00",
9716=>X"00",
9717=>X"00",
9718=>X"00",
9719=>X"00",
9720=>X"00",
9721=>X"00",
9722=>X"00",
9723=>X"00",
9724=>X"00",
9725=>X"00",
9726=>X"00",
9727=>X"00",
9728=>X"15",
9729=>X"15",
9730=>X"15",
9731=>X"15",
9732=>X"15",
9733=>X"15",
9734=>X"15",
9735=>X"15",
9736=>X"15",
9737=>X"15",
9738=>X"15",
9739=>X"15",
9740=>X"15",
9741=>X"15",
9742=>X"15",
9743=>X"15",
9744=>X"15",
9745=>X"15",
9746=>X"15",
9747=>X"15",
9748=>X"15",
9749=>X"15",
9750=>X"15",
9751=>X"15",
9752=>X"15",
9753=>X"15",
9754=>X"15",
9755=>X"15",
9756=>X"15",
9757=>X"2A",
9758=>X"2E",
9759=>X"2E",
9760=>X"2A",
9761=>X"1A",
9762=>X"1A",
9763=>X"19",
9764=>X"29",
9765=>X"19",
9766=>X"19",
9767=>X"19",
9768=>X"19",
9769=>X"19",
9770=>X"19",
9771=>X"19",
9772=>X"19",
9773=>X"19",
9774=>X"19",
9775=>X"15",
9776=>X"19",
9777=>X"19",
9778=>X"2A",
9779=>X"3E",
9780=>X"3E",
9781=>X"3E",
9782=>X"3E",
9783=>X"3E",
9784=>X"3E",
9785=>X"3E",
9786=>X"3E",
9787=>X"3E",
9788=>X"3E",
9789=>X"39",
9790=>X"2A",
9791=>X"26",
9792=>X"16",
9793=>X"16",
9794=>X"26",
9795=>X"16",
9796=>X"15",
9797=>X"15",
9798=>X"15",
9799=>X"15",
9800=>X"15",
9801=>X"15",
9802=>X"15",
9803=>X"15",
9804=>X"15",
9805=>X"15",
9806=>X"15",
9807=>X"15",
9808=>X"15",
9809=>X"15",
9810=>X"15",
9811=>X"15",
9812=>X"15",
9813=>X"15",
9814=>X"15",
9815=>X"15",
9816=>X"15",
9817=>X"15",
9818=>X"15",
9819=>X"15",
9820=>X"15",
9821=>X"15",
9822=>X"15",
9823=>X"15",
9824=>X"15",
9825=>X"15",
9826=>X"15",
9827=>X"15",
9828=>X"00",
9829=>X"00",
9830=>X"00",
9831=>X"00",
9832=>X"00",
9833=>X"00",
9834=>X"00",
9835=>X"00",
9836=>X"00",
9837=>X"00",
9838=>X"00",
9839=>X"00",
9840=>X"00",
9841=>X"00",
9842=>X"00",
9843=>X"00",
9844=>X"00",
9845=>X"00",
9846=>X"00",
9847=>X"00",
9848=>X"00",
9849=>X"00",
9850=>X"00",
9851=>X"00",
9852=>X"00",
9853=>X"00",
9854=>X"00",
9855=>X"00",
9856=>X"00",
9857=>X"00",
9858=>X"00",
9859=>X"00",
9860=>X"00",
9861=>X"00",
9862=>X"00",
9863=>X"00",
9864=>X"00",
9865=>X"00",
9866=>X"00",
9867=>X"00",
9868=>X"00",
9869=>X"00",
9870=>X"00",
9871=>X"00",
9872=>X"00",
9873=>X"00",
9874=>X"00",
9875=>X"00",
9876=>X"00",
9877=>X"00",
9878=>X"00",
9879=>X"00",
9880=>X"00",
9881=>X"00",
9882=>X"00",
9883=>X"00",
9884=>X"00",
9885=>X"00",
9886=>X"00",
9887=>X"00",
9888=>X"00",
9889=>X"00",
9890=>X"00",
9891=>X"00",
9892=>X"00",
9893=>X"00",
9894=>X"00",
9895=>X"00",
9896=>X"00",
9897=>X"00",
9898=>X"00",
9899=>X"00",
9900=>X"00",
9901=>X"00",
9902=>X"00",
9903=>X"00",
9904=>X"00",
9905=>X"00",
9906=>X"00",
9907=>X"00",
9908=>X"00",
9909=>X"00",
9910=>X"00",
9911=>X"00",
9912=>X"00",
9913=>X"00",
9914=>X"00",
9915=>X"00",
9916=>X"00",
9917=>X"00",
9918=>X"00",
9919=>X"00",
9920=>X"00",
9921=>X"00",
9922=>X"00",
9923=>X"00",
9924=>X"00",
9925=>X"00",
9926=>X"00",
9927=>X"00",
9928=>X"00",
9929=>X"00",
9930=>X"00",
9931=>X"00",
9932=>X"00",
9933=>X"00",
9934=>X"00",
9935=>X"00",
9936=>X"00",
9937=>X"00",
9938=>X"00",
9939=>X"00",
9940=>X"00",
9941=>X"00",
9942=>X"00",
9943=>X"00",
9944=>X"00",
9945=>X"00",
9946=>X"00",
9947=>X"00",
9948=>X"00",
9949=>X"00",
9950=>X"00",
9951=>X"00",
9952=>X"00",
9953=>X"00",
9954=>X"00",
9955=>X"00",
9956=>X"00",
9957=>X"00",
9958=>X"00",
9959=>X"00",
9960=>X"00",
9961=>X"00",
9962=>X"00",
9963=>X"00",
9964=>X"00",
9965=>X"00",
9966=>X"00",
9967=>X"00",
9968=>X"00",
9969=>X"00",
9970=>X"00",
9971=>X"00",
9972=>X"00",
9973=>X"00",
9974=>X"00",
9975=>X"00",
9976=>X"00",
9977=>X"00",
9978=>X"00",
9979=>X"00",
9980=>X"00",
9981=>X"00",
9982=>X"00",
9983=>X"00",
9984=>X"15",
9985=>X"15",
9986=>X"15",
9987=>X"15",
9988=>X"15",
9989=>X"15",
9990=>X"15",
9991=>X"15",
9992=>X"15",
9993=>X"15",
9994=>X"15",
9995=>X"15",
9996=>X"15",
9997=>X"15",
9998=>X"15",
9999=>X"15",
10000=>X"15",
10001=>X"15",
10002=>X"15",
10003=>X"15",
10004=>X"15",
10005=>X"15",
10006=>X"15",
10007=>X"15",
10008=>X"15",
10009=>X"15",
10010=>X"15",
10011=>X"15",
10012=>X"2A",
10013=>X"2E",
10014=>X"2E",
10015=>X"2A",
10016=>X"2A",
10017=>X"2A",
10018=>X"2A",
10019=>X"2A",
10020=>X"29",
10021=>X"19",
10022=>X"19",
10023=>X"19",
10024=>X"19",
10025=>X"19",
10026=>X"19",
10027=>X"19",
10028=>X"19",
10029=>X"19",
10030=>X"19",
10031=>X"19",
10032=>X"19",
10033=>X"29",
10034=>X"3E",
10035=>X"3E",
10036=>X"3E",
10037=>X"3E",
10038=>X"3E",
10039=>X"3E",
10040=>X"3D",
10041=>X"3D",
10042=>X"3E",
10043=>X"3E",
10044=>X"3E",
10045=>X"39",
10046=>X"39",
10047=>X"2A",
10048=>X"16",
10049=>X"16",
10050=>X"26",
10051=>X"15",
10052=>X"15",
10053=>X"15",
10054=>X"15",
10055=>X"15",
10056=>X"15",
10057=>X"15",
10058=>X"15",
10059=>X"15",
10060=>X"15",
10061=>X"15",
10062=>X"15",
10063=>X"15",
10064=>X"15",
10065=>X"15",
10066=>X"15",
10067=>X"15",
10068=>X"15",
10069=>X"15",
10070=>X"15",
10071=>X"15",
10072=>X"15",
10073=>X"15",
10074=>X"15",
10075=>X"15",
10076=>X"15",
10077=>X"15",
10078=>X"15",
10079=>X"15",
10080=>X"15",
10081=>X"15",
10082=>X"15",
10083=>X"15",
10084=>X"00",
10085=>X"00",
10086=>X"00",
10087=>X"00",
10088=>X"00",
10089=>X"00",
10090=>X"00",
10091=>X"00",
10092=>X"00",
10093=>X"00",
10094=>X"00",
10095=>X"00",
10096=>X"00",
10097=>X"00",
10098=>X"00",
10099=>X"00",
10100=>X"00",
10101=>X"00",
10102=>X"00",
10103=>X"00",
10104=>X"00",
10105=>X"00",
10106=>X"00",
10107=>X"00",
10108=>X"00",
10109=>X"00",
10110=>X"00",
10111=>X"00",
10112=>X"00",
10113=>X"00",
10114=>X"00",
10115=>X"00",
10116=>X"00",
10117=>X"00",
10118=>X"00",
10119=>X"00",
10120=>X"00",
10121=>X"00",
10122=>X"00",
10123=>X"00",
10124=>X"00",
10125=>X"00",
10126=>X"00",
10127=>X"00",
10128=>X"00",
10129=>X"00",
10130=>X"00",
10131=>X"00",
10132=>X"00",
10133=>X"00",
10134=>X"00",
10135=>X"00",
10136=>X"00",
10137=>X"00",
10138=>X"00",
10139=>X"00",
10140=>X"00",
10141=>X"00",
10142=>X"00",
10143=>X"00",
10144=>X"00",
10145=>X"00",
10146=>X"00",
10147=>X"00",
10148=>X"00",
10149=>X"00",
10150=>X"00",
10151=>X"00",
10152=>X"00",
10153=>X"00",
10154=>X"00",
10155=>X"00",
10156=>X"00",
10157=>X"00",
10158=>X"00",
10159=>X"00",
10160=>X"00",
10161=>X"00",
10162=>X"00",
10163=>X"00",
10164=>X"00",
10165=>X"00",
10166=>X"00",
10167=>X"00",
10168=>X"00",
10169=>X"00",
10170=>X"00",
10171=>X"00",
10172=>X"00",
10173=>X"00",
10174=>X"00",
10175=>X"00",
10176=>X"00",
10177=>X"00",
10178=>X"00",
10179=>X"00",
10180=>X"00",
10181=>X"00",
10182=>X"00",
10183=>X"00",
10184=>X"00",
10185=>X"00",
10186=>X"00",
10187=>X"00",
10188=>X"00",
10189=>X"00",
10190=>X"00",
10191=>X"00",
10192=>X"00",
10193=>X"00",
10194=>X"00",
10195=>X"00",
10196=>X"00",
10197=>X"00",
10198=>X"00",
10199=>X"00",
10200=>X"00",
10201=>X"00",
10202=>X"00",
10203=>X"00",
10204=>X"00",
10205=>X"00",
10206=>X"00",
10207=>X"00",
10208=>X"00",
10209=>X"00",
10210=>X"00",
10211=>X"00",
10212=>X"00",
10213=>X"00",
10214=>X"00",
10215=>X"00",
10216=>X"00",
10217=>X"00",
10218=>X"00",
10219=>X"00",
10220=>X"00",
10221=>X"00",
10222=>X"00",
10223=>X"00",
10224=>X"00",
10225=>X"00",
10226=>X"00",
10227=>X"00",
10228=>X"00",
10229=>X"00",
10230=>X"00",
10231=>X"00",
10232=>X"00",
10233=>X"00",
10234=>X"00",
10235=>X"00",
10236=>X"00",
10237=>X"00",
10238=>X"00",
10239=>X"00",
10240=>X"15",
10241=>X"15",
10242=>X"15",
10243=>X"15",
10244=>X"15",
10245=>X"15",
10246=>X"15",
10247=>X"15",
10248=>X"15",
10249=>X"15",
10250=>X"15",
10251=>X"15",
10252=>X"15",
10253=>X"15",
10254=>X"15",
10255=>X"15",
10256=>X"15",
10257=>X"15",
10258=>X"15",
10259=>X"15",
10260=>X"15",
10261=>X"15",
10262=>X"15",
10263=>X"15",
10264=>X"15",
10265=>X"15",
10266=>X"15",
10267=>X"19",
10268=>X"2E",
10269=>X"2E",
10270=>X"1A",
10271=>X"2A",
10272=>X"2A",
10273=>X"29",
10274=>X"29",
10275=>X"2A",
10276=>X"19",
10277=>X"15",
10278=>X"15",
10279=>X"15",
10280=>X"19",
10281=>X"15",
10282=>X"15",
10283=>X"19",
10284=>X"15",
10285=>X"19",
10286=>X"19",
10287=>X"19",
10288=>X"29",
10289=>X"29",
10290=>X"3E",
10291=>X"3E",
10292=>X"3E",
10293=>X"3A",
10294=>X"39",
10295=>X"39",
10296=>X"39",
10297=>X"39",
10298=>X"3D",
10299=>X"3E",
10300=>X"3E",
10301=>X"3D",
10302=>X"39",
10303=>X"29",
10304=>X"16",
10305=>X"16",
10306=>X"15",
10307=>X"15",
10308=>X"15",
10309=>X"15",
10310=>X"15",
10311=>X"15",
10312=>X"15",
10313=>X"15",
10314=>X"15",
10315=>X"15",
10316=>X"15",
10317=>X"15",
10318=>X"15",
10319=>X"15",
10320=>X"15",
10321=>X"15",
10322=>X"15",
10323=>X"15",
10324=>X"15",
10325=>X"15",
10326=>X"15",
10327=>X"15",
10328=>X"15",
10329=>X"15",
10330=>X"15",
10331=>X"15",
10332=>X"15",
10333=>X"15",
10334=>X"15",
10335=>X"15",
10336=>X"15",
10337=>X"15",
10338=>X"15",
10339=>X"15",
10340=>X"00",
10341=>X"00",
10342=>X"00",
10343=>X"00",
10344=>X"00",
10345=>X"00",
10346=>X"00",
10347=>X"00",
10348=>X"00",
10349=>X"00",
10350=>X"00",
10351=>X"00",
10352=>X"00",
10353=>X"00",
10354=>X"00",
10355=>X"00",
10356=>X"00",
10357=>X"00",
10358=>X"00",
10359=>X"00",
10360=>X"00",
10361=>X"00",
10362=>X"00",
10363=>X"00",
10364=>X"00",
10365=>X"00",
10366=>X"00",
10367=>X"00",
10368=>X"00",
10369=>X"00",
10370=>X"00",
10371=>X"00",
10372=>X"00",
10373=>X"00",
10374=>X"00",
10375=>X"00",
10376=>X"00",
10377=>X"00",
10378=>X"00",
10379=>X"00",
10380=>X"00",
10381=>X"00",
10382=>X"00",
10383=>X"00",
10384=>X"00",
10385=>X"00",
10386=>X"00",
10387=>X"00",
10388=>X"00",
10389=>X"00",
10390=>X"00",
10391=>X"00",
10392=>X"00",
10393=>X"00",
10394=>X"00",
10395=>X"00",
10396=>X"00",
10397=>X"00",
10398=>X"00",
10399=>X"00",
10400=>X"00",
10401=>X"00",
10402=>X"00",
10403=>X"00",
10404=>X"00",
10405=>X"00",
10406=>X"00",
10407=>X"00",
10408=>X"00",
10409=>X"00",
10410=>X"00",
10411=>X"00",
10412=>X"00",
10413=>X"00",
10414=>X"00",
10415=>X"00",
10416=>X"00",
10417=>X"00",
10418=>X"00",
10419=>X"00",
10420=>X"00",
10421=>X"00",
10422=>X"00",
10423=>X"00",
10424=>X"00",
10425=>X"00",
10426=>X"00",
10427=>X"00",
10428=>X"00",
10429=>X"00",
10430=>X"00",
10431=>X"00",
10432=>X"00",
10433=>X"00",
10434=>X"00",
10435=>X"00",
10436=>X"00",
10437=>X"00",
10438=>X"00",
10439=>X"00",
10440=>X"00",
10441=>X"00",
10442=>X"00",
10443=>X"00",
10444=>X"00",
10445=>X"00",
10446=>X"00",
10447=>X"00",
10448=>X"00",
10449=>X"00",
10450=>X"00",
10451=>X"00",
10452=>X"00",
10453=>X"00",
10454=>X"00",
10455=>X"00",
10456=>X"00",
10457=>X"00",
10458=>X"00",
10459=>X"00",
10460=>X"00",
10461=>X"00",
10462=>X"00",
10463=>X"00",
10464=>X"00",
10465=>X"00",
10466=>X"00",
10467=>X"00",
10468=>X"00",
10469=>X"00",
10470=>X"00",
10471=>X"00",
10472=>X"00",
10473=>X"00",
10474=>X"00",
10475=>X"00",
10476=>X"00",
10477=>X"00",
10478=>X"00",
10479=>X"00",
10480=>X"00",
10481=>X"00",
10482=>X"00",
10483=>X"00",
10484=>X"00",
10485=>X"00",
10486=>X"00",
10487=>X"00",
10488=>X"00",
10489=>X"00",
10490=>X"00",
10491=>X"00",
10492=>X"00",
10493=>X"00",
10494=>X"00",
10495=>X"00",
10496=>X"15",
10497=>X"15",
10498=>X"15",
10499=>X"15",
10500=>X"15",
10501=>X"15",
10502=>X"15",
10503=>X"15",
10504=>X"15",
10505=>X"15",
10506=>X"15",
10507=>X"15",
10508=>X"15",
10509=>X"15",
10510=>X"15",
10511=>X"15",
10512=>X"15",
10513=>X"15",
10514=>X"15",
10515=>X"15",
10516=>X"15",
10517=>X"15",
10518=>X"15",
10519=>X"15",
10520=>X"15",
10521=>X"15",
10522=>X"15",
10523=>X"1A",
10524=>X"2E",
10525=>X"2E",
10526=>X"2A",
10527=>X"29",
10528=>X"29",
10529=>X"29",
10530=>X"19",
10531=>X"15",
10532=>X"15",
10533=>X"19",
10534=>X"19",
10535=>X"15",
10536=>X"15",
10537=>X"15",
10538=>X"19",
10539=>X"15",
10540=>X"15",
10541=>X"15",
10542=>X"29",
10543=>X"29",
10544=>X"29",
10545=>X"3D",
10546=>X"3E",
10547=>X"3E",
10548=>X"3E",
10549=>X"3E",
10550=>X"3E",
10551=>X"39",
10552=>X"39",
10553=>X"39",
10554=>X"3D",
10555=>X"3D",
10556=>X"3D",
10557=>X"3D",
10558=>X"39",
10559=>X"29",
10560=>X"16",
10561=>X"16",
10562=>X"15",
10563=>X"15",
10564=>X"15",
10565=>X"15",
10566=>X"15",
10567=>X"15",
10568=>X"15",
10569=>X"15",
10570=>X"15",
10571=>X"15",
10572=>X"15",
10573=>X"15",
10574=>X"15",
10575=>X"15",
10576=>X"15",
10577=>X"15",
10578=>X"15",
10579=>X"15",
10580=>X"15",
10581=>X"15",
10582=>X"15",
10583=>X"15",
10584=>X"15",
10585=>X"15",
10586=>X"15",
10587=>X"15",
10588=>X"15",
10589=>X"15",
10590=>X"15",
10591=>X"15",
10592=>X"15",
10593=>X"15",
10594=>X"19",
10595=>X"15",
10596=>X"00",
10597=>X"00",
10598=>X"00",
10599=>X"00",
10600=>X"00",
10601=>X"00",
10602=>X"00",
10603=>X"00",
10604=>X"00",
10605=>X"00",
10606=>X"00",
10607=>X"00",
10608=>X"00",
10609=>X"00",
10610=>X"00",
10611=>X"00",
10612=>X"00",
10613=>X"00",
10614=>X"00",
10615=>X"00",
10616=>X"00",
10617=>X"00",
10618=>X"00",
10619=>X"00",
10620=>X"00",
10621=>X"00",
10622=>X"00",
10623=>X"00",
10624=>X"00",
10625=>X"00",
10626=>X"00",
10627=>X"00",
10628=>X"00",
10629=>X"00",
10630=>X"00",
10631=>X"00",
10632=>X"00",
10633=>X"00",
10634=>X"00",
10635=>X"00",
10636=>X"00",
10637=>X"00",
10638=>X"00",
10639=>X"00",
10640=>X"00",
10641=>X"00",
10642=>X"00",
10643=>X"00",
10644=>X"00",
10645=>X"00",
10646=>X"00",
10647=>X"00",
10648=>X"00",
10649=>X"00",
10650=>X"00",
10651=>X"00",
10652=>X"00",
10653=>X"00",
10654=>X"00",
10655=>X"00",
10656=>X"00",
10657=>X"00",
10658=>X"00",
10659=>X"00",
10660=>X"00",
10661=>X"00",
10662=>X"00",
10663=>X"00",
10664=>X"00",
10665=>X"00",
10666=>X"00",
10667=>X"00",
10668=>X"00",
10669=>X"00",
10670=>X"00",
10671=>X"00",
10672=>X"00",
10673=>X"00",
10674=>X"00",
10675=>X"00",
10676=>X"00",
10677=>X"00",
10678=>X"00",
10679=>X"00",
10680=>X"00",
10681=>X"00",
10682=>X"00",
10683=>X"00",
10684=>X"00",
10685=>X"00",
10686=>X"00",
10687=>X"00",
10688=>X"00",
10689=>X"00",
10690=>X"00",
10691=>X"00",
10692=>X"00",
10693=>X"00",
10694=>X"00",
10695=>X"00",
10696=>X"00",
10697=>X"00",
10698=>X"00",
10699=>X"00",
10700=>X"00",
10701=>X"00",
10702=>X"00",
10703=>X"00",
10704=>X"00",
10705=>X"00",
10706=>X"00",
10707=>X"00",
10708=>X"00",
10709=>X"00",
10710=>X"00",
10711=>X"00",
10712=>X"00",
10713=>X"00",
10714=>X"00",
10715=>X"00",
10716=>X"00",
10717=>X"00",
10718=>X"00",
10719=>X"00",
10720=>X"00",
10721=>X"00",
10722=>X"00",
10723=>X"00",
10724=>X"00",
10725=>X"00",
10726=>X"00",
10727=>X"00",
10728=>X"00",
10729=>X"00",
10730=>X"00",
10731=>X"00",
10732=>X"00",
10733=>X"00",
10734=>X"00",
10735=>X"00",
10736=>X"00",
10737=>X"00",
10738=>X"00",
10739=>X"00",
10740=>X"00",
10741=>X"00",
10742=>X"00",
10743=>X"00",
10744=>X"00",
10745=>X"00",
10746=>X"00",
10747=>X"00",
10748=>X"00",
10749=>X"00",
10750=>X"00",
10751=>X"00",
10752=>X"15",
10753=>X"15",
10754=>X"15",
10755=>X"15",
10756=>X"15",
10757=>X"15",
10758=>X"15",
10759=>X"15",
10760=>X"15",
10761=>X"15",
10762=>X"15",
10763=>X"15",
10764=>X"15",
10765=>X"15",
10766=>X"15",
10767=>X"15",
10768=>X"15",
10769=>X"15",
10770=>X"15",
10771=>X"15",
10772=>X"15",
10773=>X"15",
10774=>X"15",
10775=>X"15",
10776=>X"15",
10777=>X"15",
10778=>X"1A",
10779=>X"1A",
10780=>X"2E",
10781=>X"2A",
10782=>X"29",
10783=>X"29",
10784=>X"19",
10785=>X"19",
10786=>X"15",
10787=>X"15",
10788=>X"19",
10789=>X"19",
10790=>X"15",
10791=>X"15",
10792=>X"15",
10793=>X"15",
10794=>X"19",
10795=>X"19",
10796=>X"15",
10797=>X"15",
10798=>X"29",
10799=>X"29",
10800=>X"29",
10801=>X"3D",
10802=>X"3E",
10803=>X"3E",
10804=>X"39",
10805=>X"39",
10806=>X"39",
10807=>X"39",
10808=>X"39",
10809=>X"39",
10810=>X"3D",
10811=>X"39",
10812=>X"38",
10813=>X"3C",
10814=>X"3C",
10815=>X"39",
10816=>X"16",
10817=>X"16",
10818=>X"15",
10819=>X"15",
10820=>X"15",
10821=>X"15",
10822=>X"15",
10823=>X"15",
10824=>X"15",
10825=>X"15",
10826=>X"15",
10827=>X"15",
10828=>X"15",
10829=>X"15",
10830=>X"15",
10831=>X"15",
10832=>X"15",
10833=>X"15",
10834=>X"15",
10835=>X"15",
10836=>X"15",
10837=>X"15",
10838=>X"15",
10839=>X"15",
10840=>X"15",
10841=>X"15",
10842=>X"15",
10843=>X"15",
10844=>X"15",
10845=>X"15",
10846=>X"15",
10847=>X"15",
10848=>X"15",
10849=>X"19",
10850=>X"19",
10851=>X"19",
10852=>X"00",
10853=>X"00",
10854=>X"00",
10855=>X"00",
10856=>X"00",
10857=>X"00",
10858=>X"00",
10859=>X"00",
10860=>X"00",
10861=>X"00",
10862=>X"00",
10863=>X"00",
10864=>X"00",
10865=>X"00",
10866=>X"00",
10867=>X"00",
10868=>X"00",
10869=>X"00",
10870=>X"00",
10871=>X"00",
10872=>X"00",
10873=>X"00",
10874=>X"00",
10875=>X"00",
10876=>X"00",
10877=>X"00",
10878=>X"00",
10879=>X"00",
10880=>X"00",
10881=>X"00",
10882=>X"00",
10883=>X"00",
10884=>X"00",
10885=>X"00",
10886=>X"00",
10887=>X"00",
10888=>X"00",
10889=>X"00",
10890=>X"00",
10891=>X"00",
10892=>X"00",
10893=>X"00",
10894=>X"00",
10895=>X"00",
10896=>X"00",
10897=>X"00",
10898=>X"00",
10899=>X"00",
10900=>X"00",
10901=>X"00",
10902=>X"00",
10903=>X"00",
10904=>X"00",
10905=>X"00",
10906=>X"00",
10907=>X"00",
10908=>X"00",
10909=>X"00",
10910=>X"00",
10911=>X"00",
10912=>X"00",
10913=>X"00",
10914=>X"00",
10915=>X"00",
10916=>X"00",
10917=>X"00",
10918=>X"00",
10919=>X"00",
10920=>X"00",
10921=>X"00",
10922=>X"00",
10923=>X"00",
10924=>X"00",
10925=>X"00",
10926=>X"00",
10927=>X"00",
10928=>X"00",
10929=>X"00",
10930=>X"00",
10931=>X"00",
10932=>X"00",
10933=>X"00",
10934=>X"00",
10935=>X"00",
10936=>X"00",
10937=>X"00",
10938=>X"00",
10939=>X"00",
10940=>X"00",
10941=>X"00",
10942=>X"00",
10943=>X"00",
10944=>X"00",
10945=>X"00",
10946=>X"00",
10947=>X"00",
10948=>X"00",
10949=>X"00",
10950=>X"00",
10951=>X"00",
10952=>X"00",
10953=>X"00",
10954=>X"00",
10955=>X"00",
10956=>X"00",
10957=>X"00",
10958=>X"00",
10959=>X"00",
10960=>X"00",
10961=>X"00",
10962=>X"00",
10963=>X"00",
10964=>X"00",
10965=>X"00",
10966=>X"00",
10967=>X"00",
10968=>X"00",
10969=>X"00",
10970=>X"00",
10971=>X"00",
10972=>X"00",
10973=>X"00",
10974=>X"00",
10975=>X"00",
10976=>X"00",
10977=>X"00",
10978=>X"00",
10979=>X"00",
10980=>X"00",
10981=>X"00",
10982=>X"00",
10983=>X"00",
10984=>X"00",
10985=>X"00",
10986=>X"00",
10987=>X"00",
10988=>X"00",
10989=>X"00",
10990=>X"00",
10991=>X"00",
10992=>X"00",
10993=>X"00",
10994=>X"00",
10995=>X"00",
10996=>X"00",
10997=>X"00",
10998=>X"00",
10999=>X"00",
11000=>X"00",
11001=>X"00",
11002=>X"00",
11003=>X"00",
11004=>X"00",
11005=>X"00",
11006=>X"00",
11007=>X"00",
11008=>X"15",
11009=>X"15",
11010=>X"15",
11011=>X"15",
11012=>X"15",
11013=>X"15",
11014=>X"15",
11015=>X"15",
11016=>X"15",
11017=>X"15",
11018=>X"15",
11019=>X"15",
11020=>X"15",
11021=>X"15",
11022=>X"15",
11023=>X"15",
11024=>X"15",
11025=>X"15",
11026=>X"15",
11027=>X"15",
11028=>X"15",
11029=>X"15",
11030=>X"15",
11031=>X"15",
11032=>X"15",
11033=>X"15",
11034=>X"1A",
11035=>X"1E",
11036=>X"2E",
11037=>X"2A",
11038=>X"19",
11039=>X"19",
11040=>X"19",
11041=>X"15",
11042=>X"19",
11043=>X"29",
11044=>X"19",
11045=>X"15",
11046=>X"15",
11047=>X"15",
11048=>X"15",
11049=>X"15",
11050=>X"15",
11051=>X"15",
11052=>X"15",
11053=>X"15",
11054=>X"29",
11055=>X"29",
11056=>X"3D",
11057=>X"3D",
11058=>X"3D",
11059=>X"3D",
11060=>X"3D",
11061=>X"3D",
11062=>X"39",
11063=>X"39",
11064=>X"39",
11065=>X"39",
11066=>X"39",
11067=>X"38",
11068=>X"3C",
11069=>X"3C",
11070=>X"3C",
11071=>X"39",
11072=>X"25",
11073=>X"15",
11074=>X"15",
11075=>X"15",
11076=>X"15",
11077=>X"15",
11078=>X"15",
11079=>X"15",
11080=>X"15",
11081=>X"15",
11082=>X"15",
11083=>X"15",
11084=>X"15",
11085=>X"15",
11086=>X"15",
11087=>X"15",
11088=>X"15",
11089=>X"15",
11090=>X"15",
11091=>X"15",
11092=>X"15",
11093=>X"15",
11094=>X"15",
11095=>X"15",
11096=>X"15",
11097=>X"15",
11098=>X"15",
11099=>X"15",
11100=>X"15",
11101=>X"15",
11102=>X"19",
11103=>X"19",
11104=>X"19",
11105=>X"19",
11106=>X"19",
11107=>X"19",
11108=>X"00",
11109=>X"00",
11110=>X"00",
11111=>X"00",
11112=>X"00",
11113=>X"00",
11114=>X"00",
11115=>X"00",
11116=>X"00",
11117=>X"00",
11118=>X"00",
11119=>X"00",
11120=>X"00",
11121=>X"00",
11122=>X"00",
11123=>X"00",
11124=>X"00",
11125=>X"00",
11126=>X"00",
11127=>X"00",
11128=>X"00",
11129=>X"00",
11130=>X"00",
11131=>X"00",
11132=>X"00",
11133=>X"00",
11134=>X"00",
11135=>X"00",
11136=>X"00",
11137=>X"00",
11138=>X"00",
11139=>X"00",
11140=>X"00",
11141=>X"00",
11142=>X"00",
11143=>X"00",
11144=>X"00",
11145=>X"00",
11146=>X"00",
11147=>X"00",
11148=>X"00",
11149=>X"00",
11150=>X"00",
11151=>X"00",
11152=>X"00",
11153=>X"00",
11154=>X"00",
11155=>X"00",
11156=>X"00",
11157=>X"00",
11158=>X"00",
11159=>X"00",
11160=>X"00",
11161=>X"00",
11162=>X"00",
11163=>X"00",
11164=>X"00",
11165=>X"00",
11166=>X"00",
11167=>X"00",
11168=>X"00",
11169=>X"00",
11170=>X"00",
11171=>X"00",
11172=>X"00",
11173=>X"00",
11174=>X"00",
11175=>X"00",
11176=>X"00",
11177=>X"00",
11178=>X"00",
11179=>X"00",
11180=>X"00",
11181=>X"00",
11182=>X"00",
11183=>X"00",
11184=>X"00",
11185=>X"00",
11186=>X"00",
11187=>X"00",
11188=>X"00",
11189=>X"00",
11190=>X"00",
11191=>X"00",
11192=>X"00",
11193=>X"00",
11194=>X"00",
11195=>X"00",
11196=>X"00",
11197=>X"00",
11198=>X"00",
11199=>X"00",
11200=>X"00",
11201=>X"00",
11202=>X"00",
11203=>X"00",
11204=>X"00",
11205=>X"00",
11206=>X"00",
11207=>X"00",
11208=>X"00",
11209=>X"00",
11210=>X"00",
11211=>X"00",
11212=>X"00",
11213=>X"00",
11214=>X"00",
11215=>X"00",
11216=>X"00",
11217=>X"00",
11218=>X"00",
11219=>X"00",
11220=>X"00",
11221=>X"00",
11222=>X"00",
11223=>X"00",
11224=>X"00",
11225=>X"00",
11226=>X"00",
11227=>X"00",
11228=>X"00",
11229=>X"00",
11230=>X"00",
11231=>X"00",
11232=>X"00",
11233=>X"00",
11234=>X"00",
11235=>X"00",
11236=>X"00",
11237=>X"00",
11238=>X"00",
11239=>X"00",
11240=>X"00",
11241=>X"00",
11242=>X"00",
11243=>X"00",
11244=>X"00",
11245=>X"00",
11246=>X"00",
11247=>X"00",
11248=>X"00",
11249=>X"00",
11250=>X"00",
11251=>X"00",
11252=>X"00",
11253=>X"00",
11254=>X"00",
11255=>X"00",
11256=>X"00",
11257=>X"00",
11258=>X"00",
11259=>X"00",
11260=>X"00",
11261=>X"00",
11262=>X"00",
11263=>X"00",
11264=>X"15",
11265=>X"15",
11266=>X"15",
11267=>X"15",
11268=>X"15",
11269=>X"15",
11270=>X"15",
11271=>X"15",
11272=>X"15",
11273=>X"15",
11274=>X"15",
11275=>X"15",
11276=>X"15",
11277=>X"15",
11278=>X"15",
11279=>X"15",
11280=>X"15",
11281=>X"15",
11282=>X"15",
11283=>X"15",
11284=>X"15",
11285=>X"15",
11286=>X"15",
11287=>X"15",
11288=>X"15",
11289=>X"1A",
11290=>X"1F",
11291=>X"2E",
11292=>X"2A",
11293=>X"29",
11294=>X"19",
11295=>X"19",
11296=>X"15",
11297=>X"19",
11298=>X"19",
11299=>X"19",
11300=>X"15",
11301=>X"15",
11302=>X"15",
11303=>X"15",
11304=>X"15",
11305=>X"15",
11306=>X"15",
11307=>X"15",
11308=>X"15",
11309=>X"15",
11310=>X"29",
11311=>X"3D",
11312=>X"3E",
11313=>X"3D",
11314=>X"3D",
11315=>X"3D",
11316=>X"3D",
11317=>X"3D",
11318=>X"3D",
11319=>X"39",
11320=>X"3C",
11321=>X"38",
11322=>X"38",
11323=>X"38",
11324=>X"3C",
11325=>X"3C",
11326=>X"38",
11327=>X"39",
11328=>X"25",
11329=>X"15",
11330=>X"15",
11331=>X"15",
11332=>X"15",
11333=>X"15",
11334=>X"15",
11335=>X"15",
11336=>X"15",
11337=>X"15",
11338=>X"15",
11339=>X"15",
11340=>X"15",
11341=>X"15",
11342=>X"15",
11343=>X"15",
11344=>X"15",
11345=>X"15",
11346=>X"15",
11347=>X"15",
11348=>X"15",
11349=>X"15",
11350=>X"15",
11351=>X"15",
11352=>X"15",
11353=>X"15",
11354=>X"15",
11355=>X"19",
11356=>X"19",
11357=>X"19",
11358=>X"19",
11359=>X"19",
11360=>X"19",
11361=>X"19",
11362=>X"19",
11363=>X"19",
11364=>X"00",
11365=>X"00",
11366=>X"00",
11367=>X"00",
11368=>X"00",
11369=>X"00",
11370=>X"00",
11371=>X"00",
11372=>X"00",
11373=>X"00",
11374=>X"00",
11375=>X"00",
11376=>X"00",
11377=>X"00",
11378=>X"00",
11379=>X"00",
11380=>X"00",
11381=>X"00",
11382=>X"00",
11383=>X"00",
11384=>X"00",
11385=>X"00",
11386=>X"00",
11387=>X"00",
11388=>X"00",
11389=>X"00",
11390=>X"00",
11391=>X"00",
11392=>X"00",
11393=>X"00",
11394=>X"00",
11395=>X"00",
11396=>X"00",
11397=>X"00",
11398=>X"00",
11399=>X"00",
11400=>X"00",
11401=>X"00",
11402=>X"00",
11403=>X"00",
11404=>X"00",
11405=>X"00",
11406=>X"00",
11407=>X"00",
11408=>X"00",
11409=>X"00",
11410=>X"00",
11411=>X"00",
11412=>X"00",
11413=>X"00",
11414=>X"00",
11415=>X"00",
11416=>X"00",
11417=>X"00",
11418=>X"00",
11419=>X"00",
11420=>X"00",
11421=>X"00",
11422=>X"00",
11423=>X"00",
11424=>X"00",
11425=>X"00",
11426=>X"00",
11427=>X"00",
11428=>X"00",
11429=>X"00",
11430=>X"00",
11431=>X"00",
11432=>X"00",
11433=>X"00",
11434=>X"00",
11435=>X"00",
11436=>X"00",
11437=>X"00",
11438=>X"00",
11439=>X"00",
11440=>X"00",
11441=>X"00",
11442=>X"00",
11443=>X"00",
11444=>X"00",
11445=>X"00",
11446=>X"00",
11447=>X"00",
11448=>X"00",
11449=>X"00",
11450=>X"00",
11451=>X"00",
11452=>X"00",
11453=>X"00",
11454=>X"00",
11455=>X"00",
11456=>X"00",
11457=>X"00",
11458=>X"00",
11459=>X"00",
11460=>X"00",
11461=>X"00",
11462=>X"00",
11463=>X"00",
11464=>X"00",
11465=>X"00",
11466=>X"00",
11467=>X"00",
11468=>X"00",
11469=>X"00",
11470=>X"00",
11471=>X"00",
11472=>X"00",
11473=>X"00",
11474=>X"00",
11475=>X"00",
11476=>X"00",
11477=>X"00",
11478=>X"00",
11479=>X"00",
11480=>X"00",
11481=>X"00",
11482=>X"00",
11483=>X"00",
11484=>X"00",
11485=>X"00",
11486=>X"00",
11487=>X"00",
11488=>X"00",
11489=>X"00",
11490=>X"00",
11491=>X"00",
11492=>X"00",
11493=>X"00",
11494=>X"00",
11495=>X"00",
11496=>X"00",
11497=>X"00",
11498=>X"00",
11499=>X"00",
11500=>X"00",
11501=>X"00",
11502=>X"00",
11503=>X"00",
11504=>X"00",
11505=>X"00",
11506=>X"00",
11507=>X"00",
11508=>X"00",
11509=>X"00",
11510=>X"00",
11511=>X"00",
11512=>X"00",
11513=>X"00",
11514=>X"00",
11515=>X"00",
11516=>X"00",
11517=>X"00",
11518=>X"00",
11519=>X"00",
11520=>X"15",
11521=>X"15",
11522=>X"15",
11523=>X"15",
11524=>X"15",
11525=>X"15",
11526=>X"15",
11527=>X"15",
11528=>X"15",
11529=>X"15",
11530=>X"15",
11531=>X"15",
11532=>X"15",
11533=>X"15",
11534=>X"15",
11535=>X"15",
11536=>X"15",
11537=>X"15",
11538=>X"15",
11539=>X"15",
11540=>X"15",
11541=>X"15",
11542=>X"15",
11543=>X"15",
11544=>X"2A",
11545=>X"2F",
11546=>X"2A",
11547=>X"29",
11548=>X"29",
11549=>X"19",
11550=>X"15",
11551=>X"15",
11552=>X"15",
11553=>X"19",
11554=>X"19",
11555=>X"15",
11556=>X"15",
11557=>X"15",
11558=>X"15",
11559=>X"15",
11560=>X"15",
11561=>X"15",
11562=>X"15",
11563=>X"15",
11564=>X"15",
11565=>X"29",
11566=>X"3D",
11567=>X"3D",
11568=>X"3D",
11569=>X"3D",
11570=>X"3D",
11571=>X"3D",
11572=>X"3D",
11573=>X"3C",
11574=>X"38",
11575=>X"38",
11576=>X"3C",
11577=>X"3C",
11578=>X"38",
11579=>X"38",
11580=>X"38",
11581=>X"38",
11582=>X"3C",
11583=>X"39",
11584=>X"25",
11585=>X"15",
11586=>X"15",
11587=>X"15",
11588=>X"15",
11589=>X"15",
11590=>X"15",
11591=>X"15",
11592=>X"15",
11593=>X"15",
11594=>X"15",
11595=>X"15",
11596=>X"15",
11597=>X"15",
11598=>X"15",
11599=>X"15",
11600=>X"15",
11601=>X"15",
11602=>X"15",
11603=>X"15",
11604=>X"15",
11605=>X"15",
11606=>X"15",
11607=>X"15",
11608=>X"19",
11609=>X"15",
11610=>X"15",
11611=>X"19",
11612=>X"19",
11613=>X"19",
11614=>X"19",
11615=>X"19",
11616=>X"19",
11617=>X"19",
11618=>X"29",
11619=>X"19",
11620=>X"00",
11621=>X"00",
11622=>X"00",
11623=>X"00",
11624=>X"00",
11625=>X"00",
11626=>X"00",
11627=>X"00",
11628=>X"00",
11629=>X"00",
11630=>X"00",
11631=>X"00",
11632=>X"00",
11633=>X"00",
11634=>X"00",
11635=>X"00",
11636=>X"00",
11637=>X"00",
11638=>X"00",
11639=>X"00",
11640=>X"00",
11641=>X"00",
11642=>X"00",
11643=>X"00",
11644=>X"00",
11645=>X"00",
11646=>X"00",
11647=>X"00",
11648=>X"00",
11649=>X"00",
11650=>X"00",
11651=>X"00",
11652=>X"00",
11653=>X"00",
11654=>X"00",
11655=>X"00",
11656=>X"00",
11657=>X"00",
11658=>X"00",
11659=>X"00",
11660=>X"00",
11661=>X"00",
11662=>X"00",
11663=>X"00",
11664=>X"00",
11665=>X"00",
11666=>X"00",
11667=>X"00",
11668=>X"00",
11669=>X"00",
11670=>X"00",
11671=>X"00",
11672=>X"00",
11673=>X"00",
11674=>X"00",
11675=>X"00",
11676=>X"00",
11677=>X"00",
11678=>X"00",
11679=>X"00",
11680=>X"00",
11681=>X"00",
11682=>X"00",
11683=>X"00",
11684=>X"00",
11685=>X"00",
11686=>X"00",
11687=>X"00",
11688=>X"00",
11689=>X"00",
11690=>X"00",
11691=>X"00",
11692=>X"00",
11693=>X"00",
11694=>X"00",
11695=>X"00",
11696=>X"00",
11697=>X"00",
11698=>X"00",
11699=>X"00",
11700=>X"00",
11701=>X"00",
11702=>X"00",
11703=>X"00",
11704=>X"00",
11705=>X"00",
11706=>X"00",
11707=>X"00",
11708=>X"00",
11709=>X"00",
11710=>X"00",
11711=>X"00",
11712=>X"00",
11713=>X"00",
11714=>X"00",
11715=>X"00",
11716=>X"00",
11717=>X"00",
11718=>X"00",
11719=>X"00",
11720=>X"00",
11721=>X"00",
11722=>X"00",
11723=>X"00",
11724=>X"00",
11725=>X"00",
11726=>X"00",
11727=>X"00",
11728=>X"00",
11729=>X"00",
11730=>X"00",
11731=>X"00",
11732=>X"00",
11733=>X"00",
11734=>X"00",
11735=>X"00",
11736=>X"00",
11737=>X"00",
11738=>X"00",
11739=>X"00",
11740=>X"00",
11741=>X"00",
11742=>X"00",
11743=>X"00",
11744=>X"00",
11745=>X"00",
11746=>X"00",
11747=>X"00",
11748=>X"00",
11749=>X"00",
11750=>X"00",
11751=>X"00",
11752=>X"00",
11753=>X"00",
11754=>X"00",
11755=>X"00",
11756=>X"00",
11757=>X"00",
11758=>X"00",
11759=>X"00",
11760=>X"00",
11761=>X"00",
11762=>X"00",
11763=>X"00",
11764=>X"00",
11765=>X"00",
11766=>X"00",
11767=>X"00",
11768=>X"00",
11769=>X"00",
11770=>X"00",
11771=>X"00",
11772=>X"00",
11773=>X"00",
11774=>X"00",
11775=>X"00",
11776=>X"15",
11777=>X"15",
11778=>X"15",
11779=>X"15",
11780=>X"15",
11781=>X"15",
11782=>X"15",
11783=>X"15",
11784=>X"15",
11785=>X"15",
11786=>X"15",
11787=>X"15",
11788=>X"15",
11789=>X"15",
11790=>X"15",
11791=>X"15",
11792=>X"15",
11793=>X"15",
11794=>X"15",
11795=>X"15",
11796=>X"15",
11797=>X"15",
11798=>X"15",
11799=>X"15",
11800=>X"2A",
11801=>X"2A",
11802=>X"19",
11803=>X"19",
11804=>X"19",
11805=>X"19",
11806=>X"15",
11807=>X"19",
11808=>X"25",
11809=>X"15",
11810=>X"15",
11811=>X"15",
11812=>X"15",
11813=>X"15",
11814=>X"15",
11815=>X"15",
11816=>X"15",
11817=>X"15",
11818=>X"15",
11819=>X"15",
11820=>X"25",
11821=>X"2D",
11822=>X"3D",
11823=>X"3D",
11824=>X"3D",
11825=>X"3D",
11826=>X"3D",
11827=>X"3D",
11828=>X"38",
11829=>X"3C",
11830=>X"3C",
11831=>X"3C",
11832=>X"3C",
11833=>X"3C",
11834=>X"38",
11835=>X"38",
11836=>X"38",
11837=>X"38",
11838=>X"38",
11839=>X"38",
11840=>X"15",
11841=>X"15",
11842=>X"15",
11843=>X"15",
11844=>X"15",
11845=>X"15",
11846=>X"15",
11847=>X"15",
11848=>X"15",
11849=>X"15",
11850=>X"15",
11851=>X"15",
11852=>X"15",
11853=>X"15",
11854=>X"15",
11855=>X"15",
11856=>X"15",
11857=>X"15",
11858=>X"15",
11859=>X"15",
11860=>X"15",
11861=>X"15",
11862=>X"15",
11863=>X"15",
11864=>X"15",
11865=>X"15",
11866=>X"19",
11867=>X"19",
11868=>X"19",
11869=>X"19",
11870=>X"19",
11871=>X"19",
11872=>X"29",
11873=>X"19",
11874=>X"19",
11875=>X"19",
11876=>X"00",
11877=>X"00",
11878=>X"00",
11879=>X"00",
11880=>X"00",
11881=>X"00",
11882=>X"00",
11883=>X"00",
11884=>X"00",
11885=>X"00",
11886=>X"00",
11887=>X"00",
11888=>X"00",
11889=>X"00",
11890=>X"00",
11891=>X"00",
11892=>X"00",
11893=>X"00",
11894=>X"00",
11895=>X"00",
11896=>X"00",
11897=>X"00",
11898=>X"00",
11899=>X"00",
11900=>X"00",
11901=>X"00",
11902=>X"00",
11903=>X"00",
11904=>X"00",
11905=>X"00",
11906=>X"00",
11907=>X"00",
11908=>X"00",
11909=>X"00",
11910=>X"00",
11911=>X"00",
11912=>X"00",
11913=>X"00",
11914=>X"00",
11915=>X"00",
11916=>X"00",
11917=>X"00",
11918=>X"00",
11919=>X"00",
11920=>X"00",
11921=>X"00",
11922=>X"00",
11923=>X"00",
11924=>X"00",
11925=>X"00",
11926=>X"00",
11927=>X"00",
11928=>X"00",
11929=>X"00",
11930=>X"00",
11931=>X"00",
11932=>X"00",
11933=>X"00",
11934=>X"00",
11935=>X"00",
11936=>X"00",
11937=>X"00",
11938=>X"00",
11939=>X"00",
11940=>X"00",
11941=>X"00",
11942=>X"00",
11943=>X"00",
11944=>X"00",
11945=>X"00",
11946=>X"00",
11947=>X"00",
11948=>X"00",
11949=>X"00",
11950=>X"00",
11951=>X"00",
11952=>X"00",
11953=>X"00",
11954=>X"00",
11955=>X"00",
11956=>X"00",
11957=>X"00",
11958=>X"00",
11959=>X"00",
11960=>X"00",
11961=>X"00",
11962=>X"00",
11963=>X"00",
11964=>X"00",
11965=>X"00",
11966=>X"00",
11967=>X"00",
11968=>X"00",
11969=>X"00",
11970=>X"00",
11971=>X"00",
11972=>X"00",
11973=>X"00",
11974=>X"00",
11975=>X"00",
11976=>X"00",
11977=>X"00",
11978=>X"00",
11979=>X"00",
11980=>X"00",
11981=>X"00",
11982=>X"00",
11983=>X"00",
11984=>X"00",
11985=>X"00",
11986=>X"00",
11987=>X"00",
11988=>X"00",
11989=>X"00",
11990=>X"00",
11991=>X"00",
11992=>X"00",
11993=>X"00",
11994=>X"00",
11995=>X"00",
11996=>X"00",
11997=>X"00",
11998=>X"00",
11999=>X"00",
12000=>X"00",
12001=>X"00",
12002=>X"00",
12003=>X"00",
12004=>X"00",
12005=>X"00",
12006=>X"00",
12007=>X"00",
12008=>X"00",
12009=>X"00",
12010=>X"00",
12011=>X"00",
12012=>X"00",
12013=>X"00",
12014=>X"00",
12015=>X"00",
12016=>X"00",
12017=>X"00",
12018=>X"00",
12019=>X"00",
12020=>X"00",
12021=>X"00",
12022=>X"00",
12023=>X"00",
12024=>X"00",
12025=>X"00",
12026=>X"00",
12027=>X"00",
12028=>X"00",
12029=>X"00",
12030=>X"00",
12031=>X"00",
12032=>X"15",
12033=>X"15",
12034=>X"15",
12035=>X"15",
12036=>X"15",
12037=>X"15",
12038=>X"15",
12039=>X"15",
12040=>X"15",
12041=>X"15",
12042=>X"15",
12043=>X"15",
12044=>X"15",
12045=>X"15",
12046=>X"15",
12047=>X"15",
12048=>X"15",
12049=>X"15",
12050=>X"15",
12051=>X"15",
12052=>X"15",
12053=>X"15",
12054=>X"15",
12055=>X"15",
12056=>X"2A",
12057=>X"2A",
12058=>X"19",
12059=>X"19",
12060=>X"15",
12061=>X"15",
12062=>X"15",
12063=>X"15",
12064=>X"15",
12065=>X"15",
12066=>X"15",
12067=>X"15",
12068=>X"15",
12069=>X"15",
12070=>X"15",
12071=>X"15",
12072=>X"15",
12073=>X"15",
12074=>X"29",
12075=>X"29",
12076=>X"39",
12077=>X"3D",
12078=>X"3D",
12079=>X"3D",
12080=>X"3D",
12081=>X"3D",
12082=>X"3D",
12083=>X"3C",
12084=>X"3C",
12085=>X"3C",
12086=>X"3C",
12087=>X"3C",
12088=>X"38",
12089=>X"38",
12090=>X"38",
12091=>X"38",
12092=>X"38",
12093=>X"38",
12094=>X"38",
12095=>X"38",
12096=>X"15",
12097=>X"15",
12098=>X"15",
12099=>X"15",
12100=>X"15",
12101=>X"15",
12102=>X"15",
12103=>X"15",
12104=>X"15",
12105=>X"15",
12106=>X"15",
12107=>X"15",
12108=>X"15",
12109=>X"15",
12110=>X"15",
12111=>X"15",
12112=>X"15",
12113=>X"15",
12114=>X"15",
12115=>X"15",
12116=>X"15",
12117=>X"15",
12118=>X"19",
12119=>X"19",
12120=>X"19",
12121=>X"19",
12122=>X"19",
12123=>X"19",
12124=>X"19",
12125=>X"19",
12126=>X"19",
12127=>X"19",
12128=>X"19",
12129=>X"15",
12130=>X"29",
12131=>X"29",
12132=>X"00",
12133=>X"00",
12134=>X"00",
12135=>X"00",
12136=>X"00",
12137=>X"00",
12138=>X"00",
12139=>X"00",
12140=>X"00",
12141=>X"00",
12142=>X"00",
12143=>X"00",
12144=>X"00",
12145=>X"00",
12146=>X"00",
12147=>X"00",
12148=>X"00",
12149=>X"00",
12150=>X"00",
12151=>X"00",
12152=>X"00",
12153=>X"00",
12154=>X"00",
12155=>X"00",
12156=>X"00",
12157=>X"00",
12158=>X"00",
12159=>X"00",
12160=>X"00",
12161=>X"00",
12162=>X"00",
12163=>X"00",
12164=>X"00",
12165=>X"00",
12166=>X"00",
12167=>X"00",
12168=>X"00",
12169=>X"00",
12170=>X"00",
12171=>X"00",
12172=>X"00",
12173=>X"00",
12174=>X"00",
12175=>X"00",
12176=>X"00",
12177=>X"00",
12178=>X"00",
12179=>X"00",
12180=>X"00",
12181=>X"00",
12182=>X"00",
12183=>X"00",
12184=>X"00",
12185=>X"00",
12186=>X"00",
12187=>X"00",
12188=>X"00",
12189=>X"00",
12190=>X"00",
12191=>X"00",
12192=>X"00",
12193=>X"00",
12194=>X"00",
12195=>X"00",
12196=>X"00",
12197=>X"00",
12198=>X"00",
12199=>X"00",
12200=>X"00",
12201=>X"00",
12202=>X"00",
12203=>X"00",
12204=>X"00",
12205=>X"00",
12206=>X"00",
12207=>X"00",
12208=>X"00",
12209=>X"00",
12210=>X"00",
12211=>X"00",
12212=>X"00",
12213=>X"00",
12214=>X"00",
12215=>X"00",
12216=>X"00",
12217=>X"00",
12218=>X"00",
12219=>X"00",
12220=>X"00",
12221=>X"00",
12222=>X"00",
12223=>X"00",
12224=>X"00",
12225=>X"00",
12226=>X"00",
12227=>X"00",
12228=>X"00",
12229=>X"00",
12230=>X"00",
12231=>X"00",
12232=>X"00",
12233=>X"00",
12234=>X"00",
12235=>X"00",
12236=>X"00",
12237=>X"00",
12238=>X"00",
12239=>X"00",
12240=>X"00",
12241=>X"00",
12242=>X"00",
12243=>X"00",
12244=>X"00",
12245=>X"00",
12246=>X"00",
12247=>X"00",
12248=>X"00",
12249=>X"00",
12250=>X"00",
12251=>X"00",
12252=>X"00",
12253=>X"00",
12254=>X"00",
12255=>X"00",
12256=>X"00",
12257=>X"00",
12258=>X"00",
12259=>X"00",
12260=>X"00",
12261=>X"00",
12262=>X"00",
12263=>X"00",
12264=>X"00",
12265=>X"00",
12266=>X"00",
12267=>X"00",
12268=>X"00",
12269=>X"00",
12270=>X"00",
12271=>X"00",
12272=>X"00",
12273=>X"00",
12274=>X"00",
12275=>X"00",
12276=>X"00",
12277=>X"00",
12278=>X"00",
12279=>X"00",
12280=>X"00",
12281=>X"00",
12282=>X"00",
12283=>X"00",
12284=>X"00",
12285=>X"00",
12286=>X"00",
12287=>X"00",
12288=>X"15",
12289=>X"15",
12290=>X"15",
12291=>X"15",
12292=>X"15",
12293=>X"15",
12294=>X"15",
12295=>X"15",
12296=>X"15",
12297=>X"15",
12298=>X"15",
12299=>X"15",
12300=>X"15",
12301=>X"15",
12302=>X"15",
12303=>X"15",
12304=>X"15",
12305=>X"15",
12306=>X"15",
12307=>X"15",
12308=>X"15",
12309=>X"15",
12310=>X"15",
12311=>X"2A",
12312=>X"2A",
12313=>X"29",
12314=>X"19",
12315=>X"15",
12316=>X"15",
12317=>X"15",
12318=>X"15",
12319=>X"15",
12320=>X"15",
12321=>X"15",
12322=>X"15",
12323=>X"15",
12324=>X"15",
12325=>X"15",
12326=>X"15",
12327=>X"15",
12328=>X"15",
12329=>X"28",
12330=>X"28",
12331=>X"3D",
12332=>X"3D",
12333=>X"3D",
12334=>X"3D",
12335=>X"39",
12336=>X"3D",
12337=>X"3D",
12338=>X"38",
12339=>X"3C",
12340=>X"3C",
12341=>X"3C",
12342=>X"38",
12343=>X"38",
12344=>X"38",
12345=>X"38",
12346=>X"38",
12347=>X"38",
12348=>X"38",
12349=>X"38",
12350=>X"39",
12351=>X"29",
12352=>X"15",
12353=>X"15",
12354=>X"15",
12355=>X"15",
12356=>X"15",
12357=>X"15",
12358=>X"15",
12359=>X"15",
12360=>X"15",
12361=>X"15",
12362=>X"15",
12363=>X"15",
12364=>X"15",
12365=>X"15",
12366=>X"15",
12367=>X"15",
12368=>X"15",
12369=>X"15",
12370=>X"15",
12371=>X"15",
12372=>X"15",
12373=>X"19",
12374=>X"19",
12375=>X"19",
12376=>X"19",
12377=>X"19",
12378=>X"29",
12379=>X"19",
12380=>X"29",
12381=>X"19",
12382=>X"19",
12383=>X"19",
12384=>X"19",
12385=>X"19",
12386=>X"29",
12387=>X"29",
12388=>X"00",
12389=>X"00",
12390=>X"00",
12391=>X"00",
12392=>X"00",
12393=>X"00",
12394=>X"00",
12395=>X"00",
12396=>X"00",
12397=>X"00",
12398=>X"00",
12399=>X"00",
12400=>X"00",
12401=>X"00",
12402=>X"00",
12403=>X"00",
12404=>X"00",
12405=>X"00",
12406=>X"00",
12407=>X"00",
12408=>X"00",
12409=>X"00",
12410=>X"00",
12411=>X"00",
12412=>X"00",
12413=>X"00",
12414=>X"00",
12415=>X"00",
12416=>X"00",
12417=>X"00",
12418=>X"00",
12419=>X"00",
12420=>X"00",
12421=>X"00",
12422=>X"00",
12423=>X"00",
12424=>X"00",
12425=>X"00",
12426=>X"00",
12427=>X"00",
12428=>X"00",
12429=>X"00",
12430=>X"00",
12431=>X"00",
12432=>X"00",
12433=>X"00",
12434=>X"00",
12435=>X"00",
12436=>X"00",
12437=>X"00",
12438=>X"00",
12439=>X"00",
12440=>X"00",
12441=>X"00",
12442=>X"00",
12443=>X"00",
12444=>X"00",
12445=>X"00",
12446=>X"00",
12447=>X"00",
12448=>X"00",
12449=>X"00",
12450=>X"00",
12451=>X"00",
12452=>X"00",
12453=>X"00",
12454=>X"00",
12455=>X"00",
12456=>X"00",
12457=>X"00",
12458=>X"00",
12459=>X"00",
12460=>X"00",
12461=>X"00",
12462=>X"00",
12463=>X"00",
12464=>X"00",
12465=>X"00",
12466=>X"00",
12467=>X"00",
12468=>X"00",
12469=>X"00",
12470=>X"00",
12471=>X"00",
12472=>X"00",
12473=>X"00",
12474=>X"00",
12475=>X"00",
12476=>X"00",
12477=>X"00",
12478=>X"00",
12479=>X"00",
12480=>X"00",
12481=>X"00",
12482=>X"00",
12483=>X"00",
12484=>X"00",
12485=>X"00",
12486=>X"00",
12487=>X"00",
12488=>X"00",
12489=>X"00",
12490=>X"00",
12491=>X"00",
12492=>X"00",
12493=>X"00",
12494=>X"00",
12495=>X"00",
12496=>X"00",
12497=>X"00",
12498=>X"00",
12499=>X"00",
12500=>X"00",
12501=>X"00",
12502=>X"00",
12503=>X"00",
12504=>X"00",
12505=>X"00",
12506=>X"00",
12507=>X"00",
12508=>X"00",
12509=>X"00",
12510=>X"00",
12511=>X"00",
12512=>X"00",
12513=>X"00",
12514=>X"00",
12515=>X"00",
12516=>X"00",
12517=>X"00",
12518=>X"00",
12519=>X"00",
12520=>X"00",
12521=>X"00",
12522=>X"00",
12523=>X"00",
12524=>X"00",
12525=>X"00",
12526=>X"00",
12527=>X"00",
12528=>X"00",
12529=>X"00",
12530=>X"00",
12531=>X"00",
12532=>X"00",
12533=>X"00",
12534=>X"00",
12535=>X"00",
12536=>X"00",
12537=>X"00",
12538=>X"00",
12539=>X"00",
12540=>X"00",
12541=>X"00",
12542=>X"00",
12543=>X"00",
12544=>X"15",
12545=>X"15",
12546=>X"15",
12547=>X"15",
12548=>X"15",
12549=>X"15",
12550=>X"15",
12551=>X"15",
12552=>X"15",
12553=>X"15",
12554=>X"15",
12555=>X"15",
12556=>X"15",
12557=>X"15",
12558=>X"15",
12559=>X"15",
12560=>X"15",
12561=>X"15",
12562=>X"15",
12563=>X"15",
12564=>X"15",
12565=>X"25",
12566=>X"19",
12567=>X"19",
12568=>X"15",
12569=>X"15",
12570=>X"15",
12571=>X"15",
12572=>X"15",
12573=>X"15",
12574=>X"15",
12575=>X"15",
12576=>X"15",
12577=>X"15",
12578=>X"15",
12579=>X"15",
12580=>X"15",
12581=>X"15",
12582=>X"15",
12583=>X"29",
12584=>X"29",
12585=>X"2C",
12586=>X"3C",
12587=>X"3C",
12588=>X"38",
12589=>X"3D",
12590=>X"3D",
12591=>X"3D",
12592=>X"39",
12593=>X"3C",
12594=>X"38",
12595=>X"38",
12596=>X"38",
12597=>X"38",
12598=>X"38",
12599=>X"38",
12600=>X"38",
12601=>X"38",
12602=>X"38",
12603=>X"38",
12604=>X"38",
12605=>X"38",
12606=>X"39",
12607=>X"29",
12608=>X"15",
12609=>X"15",
12610=>X"15",
12611=>X"15",
12612=>X"15",
12613=>X"15",
12614=>X"15",
12615=>X"15",
12616=>X"15",
12617=>X"15",
12618=>X"15",
12619=>X"15",
12620=>X"15",
12621=>X"15",
12622=>X"15",
12623=>X"15",
12624=>X"15",
12625=>X"15",
12626=>X"15",
12627=>X"15",
12628=>X"15",
12629=>X"15",
12630=>X"19",
12631=>X"29",
12632=>X"19",
12633=>X"19",
12634=>X"19",
12635=>X"19",
12636=>X"19",
12637=>X"19",
12638=>X"29",
12639=>X"19",
12640=>X"19",
12641=>X"19",
12642=>X"19",
12643=>X"19",
12644=>X"00",
12645=>X"00",
12646=>X"00",
12647=>X"00",
12648=>X"00",
12649=>X"00",
12650=>X"00",
12651=>X"00",
12652=>X"00",
12653=>X"00",
12654=>X"00",
12655=>X"00",
12656=>X"00",
12657=>X"00",
12658=>X"00",
12659=>X"00",
12660=>X"00",
12661=>X"00",
12662=>X"00",
12663=>X"00",
12664=>X"00",
12665=>X"00",
12666=>X"00",
12667=>X"00",
12668=>X"00",
12669=>X"00",
12670=>X"00",
12671=>X"00",
12672=>X"00",
12673=>X"00",
12674=>X"00",
12675=>X"00",
12676=>X"00",
12677=>X"00",
12678=>X"00",
12679=>X"00",
12680=>X"00",
12681=>X"00",
12682=>X"00",
12683=>X"00",
12684=>X"00",
12685=>X"00",
12686=>X"00",
12687=>X"00",
12688=>X"00",
12689=>X"00",
12690=>X"00",
12691=>X"00",
12692=>X"00",
12693=>X"00",
12694=>X"00",
12695=>X"00",
12696=>X"00",
12697=>X"00",
12698=>X"00",
12699=>X"00",
12700=>X"00",
12701=>X"00",
12702=>X"00",
12703=>X"00",
12704=>X"00",
12705=>X"00",
12706=>X"00",
12707=>X"00",
12708=>X"00",
12709=>X"00",
12710=>X"00",
12711=>X"00",
12712=>X"00",
12713=>X"00",
12714=>X"00",
12715=>X"00",
12716=>X"00",
12717=>X"00",
12718=>X"00",
12719=>X"00",
12720=>X"00",
12721=>X"00",
12722=>X"00",
12723=>X"00",
12724=>X"00",
12725=>X"00",
12726=>X"00",
12727=>X"00",
12728=>X"00",
12729=>X"00",
12730=>X"00",
12731=>X"00",
12732=>X"00",
12733=>X"00",
12734=>X"00",
12735=>X"00",
12736=>X"00",
12737=>X"00",
12738=>X"00",
12739=>X"00",
12740=>X"00",
12741=>X"00",
12742=>X"00",
12743=>X"00",
12744=>X"00",
12745=>X"00",
12746=>X"00",
12747=>X"00",
12748=>X"00",
12749=>X"00",
12750=>X"00",
12751=>X"00",
12752=>X"00",
12753=>X"00",
12754=>X"00",
12755=>X"00",
12756=>X"00",
12757=>X"00",
12758=>X"00",
12759=>X"00",
12760=>X"00",
12761=>X"00",
12762=>X"00",
12763=>X"00",
12764=>X"00",
12765=>X"00",
12766=>X"00",
12767=>X"00",
12768=>X"00",
12769=>X"00",
12770=>X"00",
12771=>X"00",
12772=>X"00",
12773=>X"00",
12774=>X"00",
12775=>X"00",
12776=>X"00",
12777=>X"00",
12778=>X"00",
12779=>X"00",
12780=>X"00",
12781=>X"00",
12782=>X"00",
12783=>X"00",
12784=>X"00",
12785=>X"00",
12786=>X"00",
12787=>X"00",
12788=>X"00",
12789=>X"00",
12790=>X"00",
12791=>X"00",
12792=>X"00",
12793=>X"00",
12794=>X"00",
12795=>X"00",
12796=>X"00",
12797=>X"00",
12798=>X"00",
12799=>X"00",
12800=>X"15",
12801=>X"15",
12802=>X"15",
12803=>X"15",
12804=>X"15",
12805=>X"15",
12806=>X"15",
12807=>X"15",
12808=>X"15",
12809=>X"15",
12810=>X"15",
12811=>X"15",
12812=>X"15",
12813=>X"15",
12814=>X"15",
12815=>X"15",
12816=>X"15",
12817=>X"15",
12818=>X"15",
12819=>X"15",
12820=>X"29",
12821=>X"25",
12822=>X"19",
12823=>X"15",
12824=>X"15",
12825=>X"15",
12826=>X"15",
12827=>X"15",
12828=>X"15",
12829=>X"15",
12830=>X"15",
12831=>X"15",
12832=>X"15",
12833=>X"15",
12834=>X"16",
12835=>X"16",
12836=>X"16",
12837=>X"19",
12838=>X"29",
12839=>X"29",
12840=>X"3D",
12841=>X"3D",
12842=>X"3C",
12843=>X"38",
12844=>X"3C",
12845=>X"3C",
12846=>X"3C",
12847=>X"3C",
12848=>X"38",
12849=>X"38",
12850=>X"38",
12851=>X"38",
12852=>X"38",
12853=>X"38",
12854=>X"38",
12855=>X"38",
12856=>X"38",
12857=>X"38",
12858=>X"38",
12859=>X"38",
12860=>X"38",
12861=>X"38",
12862=>X"29",
12863=>X"25",
12864=>X"15",
12865=>X"15",
12866=>X"15",
12867=>X"15",
12868=>X"15",
12869=>X"15",
12870=>X"15",
12871=>X"15",
12872=>X"15",
12873=>X"15",
12874=>X"15",
12875=>X"15",
12876=>X"15",
12877=>X"15",
12878=>X"15",
12879=>X"15",
12880=>X"15",
12881=>X"15",
12882=>X"19",
12883=>X"15",
12884=>X"19",
12885=>X"19",
12886=>X"19",
12887=>X"29",
12888=>X"19",
12889=>X"29",
12890=>X"19",
12891=>X"19",
12892=>X"19",
12893=>X"19",
12894=>X"29",
12895=>X"19",
12896=>X"19",
12897=>X"19",
12898=>X"19",
12899=>X"19",
12900=>X"00",
12901=>X"00",
12902=>X"00",
12903=>X"00",
12904=>X"00",
12905=>X"00",
12906=>X"00",
12907=>X"00",
12908=>X"00",
12909=>X"00",
12910=>X"00",
12911=>X"00",
12912=>X"00",
12913=>X"00",
12914=>X"00",
12915=>X"00",
12916=>X"00",
12917=>X"00",
12918=>X"00",
12919=>X"00",
12920=>X"00",
12921=>X"00",
12922=>X"00",
12923=>X"00",
12924=>X"00",
12925=>X"00",
12926=>X"00",
12927=>X"00",
12928=>X"00",
12929=>X"00",
12930=>X"00",
12931=>X"00",
12932=>X"00",
12933=>X"00",
12934=>X"00",
12935=>X"00",
12936=>X"00",
12937=>X"00",
12938=>X"00",
12939=>X"00",
12940=>X"00",
12941=>X"00",
12942=>X"00",
12943=>X"00",
12944=>X"00",
12945=>X"00",
12946=>X"00",
12947=>X"00",
12948=>X"00",
12949=>X"00",
12950=>X"00",
12951=>X"00",
12952=>X"00",
12953=>X"00",
12954=>X"00",
12955=>X"00",
12956=>X"00",
12957=>X"00",
12958=>X"00",
12959=>X"00",
12960=>X"00",
12961=>X"00",
12962=>X"00",
12963=>X"00",
12964=>X"00",
12965=>X"00",
12966=>X"00",
12967=>X"00",
12968=>X"00",
12969=>X"00",
12970=>X"00",
12971=>X"00",
12972=>X"00",
12973=>X"00",
12974=>X"00",
12975=>X"00",
12976=>X"00",
12977=>X"00",
12978=>X"00",
12979=>X"00",
12980=>X"00",
12981=>X"00",
12982=>X"00",
12983=>X"00",
12984=>X"00",
12985=>X"00",
12986=>X"00",
12987=>X"00",
12988=>X"00",
12989=>X"00",
12990=>X"00",
12991=>X"00",
12992=>X"00",
12993=>X"00",
12994=>X"00",
12995=>X"00",
12996=>X"00",
12997=>X"00",
12998=>X"00",
12999=>X"00",
13000=>X"00",
13001=>X"00",
13002=>X"00",
13003=>X"00",
13004=>X"00",
13005=>X"00",
13006=>X"00",
13007=>X"00",
13008=>X"00",
13009=>X"00",
13010=>X"00",
13011=>X"00",
13012=>X"00",
13013=>X"00",
13014=>X"00",
13015=>X"00",
13016=>X"00",
13017=>X"00",
13018=>X"00",
13019=>X"00",
13020=>X"00",
13021=>X"00",
13022=>X"00",
13023=>X"00",
13024=>X"00",
13025=>X"00",
13026=>X"00",
13027=>X"00",
13028=>X"00",
13029=>X"00",
13030=>X"00",
13031=>X"00",
13032=>X"00",
13033=>X"00",
13034=>X"00",
13035=>X"00",
13036=>X"00",
13037=>X"00",
13038=>X"00",
13039=>X"00",
13040=>X"00",
13041=>X"00",
13042=>X"00",
13043=>X"00",
13044=>X"00",
13045=>X"00",
13046=>X"00",
13047=>X"00",
13048=>X"00",
13049=>X"00",
13050=>X"00",
13051=>X"00",
13052=>X"00",
13053=>X"00",
13054=>X"00",
13055=>X"00",
13056=>X"15",
13057=>X"15",
13058=>X"15",
13059=>X"15",
13060=>X"15",
13061=>X"15",
13062=>X"15",
13063=>X"15",
13064=>X"15",
13065=>X"15",
13066=>X"15",
13067=>X"15",
13068=>X"15",
13069=>X"15",
13070=>X"15",
13071=>X"15",
13072=>X"15",
13073=>X"15",
13074=>X"15",
13075=>X"16",
13076=>X"29",
13077=>X"15",
13078=>X"15",
13079=>X"15",
13080=>X"15",
13081=>X"15",
13082=>X"16",
13083=>X"16",
13084=>X"1B",
13085=>X"1B",
13086=>X"1B",
13087=>X"1B",
13088=>X"1B",
13089=>X"1B",
13090=>X"1B",
13091=>X"1B",
13092=>X"1B",
13093=>X"1A",
13094=>X"29",
13095=>X"29",
13096=>X"3D",
13097=>X"39",
13098=>X"3C",
13099=>X"3C",
13100=>X"3C",
13101=>X"3C",
13102=>X"38",
13103=>X"3C",
13104=>X"38",
13105=>X"38",
13106=>X"38",
13107=>X"38",
13108=>X"38",
13109=>X"38",
13110=>X"38",
13111=>X"38",
13112=>X"38",
13113=>X"38",
13114=>X"38",
13115=>X"38",
13116=>X"38",
13117=>X"39",
13118=>X"25",
13119=>X"15",
13120=>X"15",
13121=>X"15",
13122=>X"15",
13123=>X"15",
13124=>X"15",
13125=>X"15",
13126=>X"15",
13127=>X"15",
13128=>X"15",
13129=>X"15",
13130=>X"15",
13131=>X"15",
13132=>X"15",
13133=>X"15",
13134=>X"15",
13135=>X"15",
13136=>X"15",
13137=>X"19",
13138=>X"19",
13139=>X"19",
13140=>X"19",
13141=>X"19",
13142=>X"29",
13143=>X"19",
13144=>X"19",
13145=>X"29",
13146=>X"19",
13147=>X"19",
13148=>X"19",
13149=>X"15",
13150=>X"19",
13151=>X"15",
13152=>X"19",
13153=>X"19",
13154=>X"19",
13155=>X"19",
13156=>X"00",
13157=>X"00",
13158=>X"00",
13159=>X"00",
13160=>X"00",
13161=>X"00",
13162=>X"00",
13163=>X"00",
13164=>X"00",
13165=>X"00",
13166=>X"00",
13167=>X"00",
13168=>X"00",
13169=>X"00",
13170=>X"00",
13171=>X"00",
13172=>X"00",
13173=>X"00",
13174=>X"00",
13175=>X"00",
13176=>X"00",
13177=>X"00",
13178=>X"00",
13179=>X"00",
13180=>X"00",
13181=>X"00",
13182=>X"00",
13183=>X"00",
13184=>X"00",
13185=>X"00",
13186=>X"00",
13187=>X"00",
13188=>X"00",
13189=>X"00",
13190=>X"00",
13191=>X"00",
13192=>X"00",
13193=>X"00",
13194=>X"00",
13195=>X"00",
13196=>X"00",
13197=>X"00",
13198=>X"00",
13199=>X"00",
13200=>X"00",
13201=>X"00",
13202=>X"00",
13203=>X"00",
13204=>X"00",
13205=>X"00",
13206=>X"00",
13207=>X"00",
13208=>X"00",
13209=>X"00",
13210=>X"00",
13211=>X"00",
13212=>X"00",
13213=>X"00",
13214=>X"00",
13215=>X"00",
13216=>X"00",
13217=>X"00",
13218=>X"00",
13219=>X"00",
13220=>X"00",
13221=>X"00",
13222=>X"00",
13223=>X"00",
13224=>X"00",
13225=>X"00",
13226=>X"00",
13227=>X"00",
13228=>X"00",
13229=>X"00",
13230=>X"00",
13231=>X"00",
13232=>X"00",
13233=>X"00",
13234=>X"00",
13235=>X"00",
13236=>X"00",
13237=>X"00",
13238=>X"00",
13239=>X"00",
13240=>X"00",
13241=>X"00",
13242=>X"00",
13243=>X"00",
13244=>X"00",
13245=>X"00",
13246=>X"00",
13247=>X"00",
13248=>X"00",
13249=>X"00",
13250=>X"00",
13251=>X"00",
13252=>X"00",
13253=>X"00",
13254=>X"00",
13255=>X"00",
13256=>X"00",
13257=>X"00",
13258=>X"00",
13259=>X"00",
13260=>X"00",
13261=>X"00",
13262=>X"00",
13263=>X"00",
13264=>X"00",
13265=>X"00",
13266=>X"00",
13267=>X"00",
13268=>X"00",
13269=>X"00",
13270=>X"00",
13271=>X"00",
13272=>X"00",
13273=>X"00",
13274=>X"00",
13275=>X"00",
13276=>X"00",
13277=>X"00",
13278=>X"00",
13279=>X"00",
13280=>X"00",
13281=>X"00",
13282=>X"00",
13283=>X"00",
13284=>X"00",
13285=>X"00",
13286=>X"00",
13287=>X"00",
13288=>X"00",
13289=>X"00",
13290=>X"00",
13291=>X"00",
13292=>X"00",
13293=>X"00",
13294=>X"00",
13295=>X"00",
13296=>X"00",
13297=>X"00",
13298=>X"00",
13299=>X"00",
13300=>X"00",
13301=>X"00",
13302=>X"00",
13303=>X"00",
13304=>X"00",
13305=>X"00",
13306=>X"00",
13307=>X"00",
13308=>X"00",
13309=>X"00",
13310=>X"00",
13311=>X"00",
13312=>X"15",
13313=>X"15",
13314=>X"15",
13315=>X"15",
13316=>X"15",
13317=>X"15",
13318=>X"15",
13319=>X"15",
13320=>X"15",
13321=>X"15",
13322=>X"15",
13323=>X"14",
13324=>X"14",
13325=>X"15",
13326=>X"14",
13327=>X"15",
13328=>X"15",
13329=>X"15",
13330=>X"15",
13331=>X"16",
13332=>X"15",
13333=>X"15",
13334=>X"15",
13335=>X"15",
13336=>X"16",
13337=>X"1A",
13338=>X"1B",
13339=>X"1B",
13340=>X"1B",
13341=>X"1B",
13342=>X"1B",
13343=>X"1B",
13344=>X"1B",
13345=>X"1B",
13346=>X"1B",
13347=>X"1B",
13348=>X"1B",
13349=>X"1A",
13350=>X"29",
13351=>X"2A",
13352=>X"3D",
13353=>X"3D",
13354=>X"3C",
13355=>X"3C",
13356=>X"38",
13357=>X"38",
13358=>X"38",
13359=>X"38",
13360=>X"38",
13361=>X"38",
13362=>X"38",
13363=>X"38",
13364=>X"38",
13365=>X"38",
13366=>X"38",
13367=>X"38",
13368=>X"38",
13369=>X"38",
13370=>X"38",
13371=>X"38",
13372=>X"39",
13373=>X"29",
13374=>X"15",
13375=>X"15",
13376=>X"15",
13377=>X"15",
13378=>X"15",
13379=>X"15",
13380=>X"15",
13381=>X"15",
13382=>X"15",
13383=>X"15",
13384=>X"15",
13385=>X"15",
13386=>X"15",
13387=>X"15",
13388=>X"15",
13389=>X"15",
13390=>X"15",
13391=>X"19",
13392=>X"19",
13393=>X"19",
13394=>X"15",
13395=>X"29",
13396=>X"19",
13397=>X"19",
13398=>X"25",
13399=>X"19",
13400=>X"19",
13401=>X"19",
13402=>X"19",
13403=>X"19",
13404=>X"19",
13405=>X"15",
13406=>X"19",
13407=>X"15",
13408=>X"19",
13409=>X"15",
13410=>X"19",
13411=>X"19",
13412=>X"00",
13413=>X"00",
13414=>X"00",
13415=>X"00",
13416=>X"00",
13417=>X"00",
13418=>X"00",
13419=>X"00",
13420=>X"00",
13421=>X"00",
13422=>X"00",
13423=>X"00",
13424=>X"00",
13425=>X"00",
13426=>X"00",
13427=>X"00",
13428=>X"00",
13429=>X"00",
13430=>X"00",
13431=>X"00",
13432=>X"00",
13433=>X"00",
13434=>X"00",
13435=>X"00",
13436=>X"00",
13437=>X"00",
13438=>X"00",
13439=>X"00",
13440=>X"00",
13441=>X"00",
13442=>X"00",
13443=>X"00",
13444=>X"00",
13445=>X"00",
13446=>X"00",
13447=>X"00",
13448=>X"00",
13449=>X"00",
13450=>X"00",
13451=>X"00",
13452=>X"00",
13453=>X"00",
13454=>X"00",
13455=>X"00",
13456=>X"00",
13457=>X"00",
13458=>X"00",
13459=>X"00",
13460=>X"00",
13461=>X"00",
13462=>X"00",
13463=>X"00",
13464=>X"00",
13465=>X"00",
13466=>X"00",
13467=>X"00",
13468=>X"00",
13469=>X"00",
13470=>X"00",
13471=>X"00",
13472=>X"00",
13473=>X"00",
13474=>X"00",
13475=>X"00",
13476=>X"00",
13477=>X"00",
13478=>X"00",
13479=>X"00",
13480=>X"00",
13481=>X"00",
13482=>X"00",
13483=>X"00",
13484=>X"00",
13485=>X"00",
13486=>X"00",
13487=>X"00",
13488=>X"00",
13489=>X"00",
13490=>X"00",
13491=>X"00",
13492=>X"00",
13493=>X"00",
13494=>X"00",
13495=>X"00",
13496=>X"00",
13497=>X"00",
13498=>X"00",
13499=>X"00",
13500=>X"00",
13501=>X"00",
13502=>X"00",
13503=>X"00",
13504=>X"00",
13505=>X"00",
13506=>X"00",
13507=>X"00",
13508=>X"00",
13509=>X"00",
13510=>X"00",
13511=>X"00",
13512=>X"00",
13513=>X"00",
13514=>X"00",
13515=>X"00",
13516=>X"00",
13517=>X"00",
13518=>X"00",
13519=>X"00",
13520=>X"00",
13521=>X"00",
13522=>X"00",
13523=>X"00",
13524=>X"00",
13525=>X"00",
13526=>X"00",
13527=>X"00",
13528=>X"00",
13529=>X"00",
13530=>X"00",
13531=>X"00",
13532=>X"00",
13533=>X"00",
13534=>X"00",
13535=>X"00",
13536=>X"00",
13537=>X"00",
13538=>X"00",
13539=>X"00",
13540=>X"00",
13541=>X"00",
13542=>X"00",
13543=>X"00",
13544=>X"00",
13545=>X"00",
13546=>X"00",
13547=>X"00",
13548=>X"00",
13549=>X"00",
13550=>X"00",
13551=>X"00",
13552=>X"00",
13553=>X"00",
13554=>X"00",
13555=>X"00",
13556=>X"00",
13557=>X"00",
13558=>X"00",
13559=>X"00",
13560=>X"00",
13561=>X"00",
13562=>X"00",
13563=>X"00",
13564=>X"00",
13565=>X"00",
13566=>X"00",
13567=>X"00",
13568=>X"15",
13569=>X"15",
13570=>X"15",
13571=>X"15",
13572=>X"15",
13573=>X"15",
13574=>X"15",
13575=>X"15",
13576=>X"15",
13577=>X"15",
13578=>X"15",
13579=>X"14",
13580=>X"14",
13581=>X"14",
13582=>X"14",
13583=>X"15",
13584=>X"15",
13585=>X"15",
13586=>X"15",
13587=>X"15",
13588=>X"15",
13589=>X"15",
13590=>X"15",
13591=>X"16",
13592=>X"1A",
13593=>X"1B",
13594=>X"1B",
13595=>X"1B",
13596=>X"1B",
13597=>X"1B",
13598=>X"1B",
13599=>X"1B",
13600=>X"1B",
13601=>X"1B",
13602=>X"1B",
13603=>X"1B",
13604=>X"1B",
13605=>X"2B",
13606=>X"3E",
13607=>X"3E",
13608=>X"3D",
13609=>X"3D",
13610=>X"38",
13611=>X"38",
13612=>X"38",
13613=>X"38",
13614=>X"38",
13615=>X"38",
13616=>X"38",
13617=>X"38",
13618=>X"38",
13619=>X"38",
13620=>X"38",
13621=>X"38",
13622=>X"38",
13623=>X"38",
13624=>X"38",
13625=>X"38",
13626=>X"38",
13627=>X"29",
13628=>X"29",
13629=>X"15",
13630=>X"15",
13631=>X"15",
13632=>X"15",
13633=>X"15",
13634=>X"15",
13635=>X"15",
13636=>X"15",
13637=>X"15",
13638=>X"15",
13639=>X"15",
13640=>X"15",
13641=>X"15",
13642=>X"15",
13643=>X"15",
13644=>X"15",
13645=>X"15",
13646=>X"15",
13647=>X"19",
13648=>X"19",
13649=>X"15",
13650=>X"19",
13651=>X"19",
13652=>X"19",
13653=>X"19",
13654=>X"15",
13655=>X"19",
13656=>X"19",
13657=>X"15",
13658=>X"19",
13659=>X"15",
13660=>X"15",
13661=>X"15",
13662=>X"15",
13663=>X"15",
13664=>X"15",
13665=>X"15",
13666=>X"15",
13667=>X"15",
13668=>X"00",
13669=>X"00",
13670=>X"00",
13671=>X"00",
13672=>X"00",
13673=>X"00",
13674=>X"00",
13675=>X"00",
13676=>X"00",
13677=>X"00",
13678=>X"00",
13679=>X"00",
13680=>X"00",
13681=>X"00",
13682=>X"00",
13683=>X"00",
13684=>X"00",
13685=>X"00",
13686=>X"00",
13687=>X"00",
13688=>X"00",
13689=>X"00",
13690=>X"00",
13691=>X"00",
13692=>X"00",
13693=>X"00",
13694=>X"00",
13695=>X"00",
13696=>X"00",
13697=>X"00",
13698=>X"00",
13699=>X"00",
13700=>X"00",
13701=>X"00",
13702=>X"00",
13703=>X"00",
13704=>X"00",
13705=>X"00",
13706=>X"00",
13707=>X"00",
13708=>X"00",
13709=>X"00",
13710=>X"00",
13711=>X"00",
13712=>X"00",
13713=>X"00",
13714=>X"00",
13715=>X"00",
13716=>X"00",
13717=>X"00",
13718=>X"00",
13719=>X"00",
13720=>X"00",
13721=>X"00",
13722=>X"00",
13723=>X"00",
13724=>X"00",
13725=>X"00",
13726=>X"00",
13727=>X"00",
13728=>X"00",
13729=>X"00",
13730=>X"00",
13731=>X"00",
13732=>X"00",
13733=>X"00",
13734=>X"00",
13735=>X"00",
13736=>X"00",
13737=>X"00",
13738=>X"00",
13739=>X"00",
13740=>X"00",
13741=>X"00",
13742=>X"00",
13743=>X"00",
13744=>X"00",
13745=>X"00",
13746=>X"00",
13747=>X"00",
13748=>X"00",
13749=>X"00",
13750=>X"00",
13751=>X"00",
13752=>X"00",
13753=>X"00",
13754=>X"00",
13755=>X"00",
13756=>X"00",
13757=>X"00",
13758=>X"00",
13759=>X"00",
13760=>X"00",
13761=>X"00",
13762=>X"00",
13763=>X"00",
13764=>X"00",
13765=>X"00",
13766=>X"00",
13767=>X"00",
13768=>X"00",
13769=>X"00",
13770=>X"00",
13771=>X"00",
13772=>X"00",
13773=>X"00",
13774=>X"00",
13775=>X"00",
13776=>X"00",
13777=>X"00",
13778=>X"00",
13779=>X"00",
13780=>X"00",
13781=>X"00",
13782=>X"00",
13783=>X"00",
13784=>X"00",
13785=>X"00",
13786=>X"00",
13787=>X"00",
13788=>X"00",
13789=>X"00",
13790=>X"00",
13791=>X"00",
13792=>X"00",
13793=>X"00",
13794=>X"00",
13795=>X"00",
13796=>X"00",
13797=>X"00",
13798=>X"00",
13799=>X"00",
13800=>X"00",
13801=>X"00",
13802=>X"00",
13803=>X"00",
13804=>X"00",
13805=>X"00",
13806=>X"00",
13807=>X"00",
13808=>X"00",
13809=>X"00",
13810=>X"00",
13811=>X"00",
13812=>X"00",
13813=>X"00",
13814=>X"00",
13815=>X"00",
13816=>X"00",
13817=>X"00",
13818=>X"00",
13819=>X"00",
13820=>X"00",
13821=>X"00",
13822=>X"00",
13823=>X"00",
13824=>X"15",
13825=>X"15",
13826=>X"15",
13827=>X"15",
13828=>X"15",
13829=>X"15",
13830=>X"15",
13831=>X"15",
13832=>X"15",
13833=>X"15",
13834=>X"14",
13835=>X"14",
13836=>X"14",
13837=>X"14",
13838=>X"14",
13839=>X"14",
13840=>X"15",
13841=>X"15",
13842=>X"15",
13843=>X"15",
13844=>X"15",
13845=>X"15",
13846=>X"05",
13847=>X"16",
13848=>X"1B",
13849=>X"1B",
13850=>X"1B",
13851=>X"1B",
13852=>X"1B",
13853=>X"1B",
13854=>X"1B",
13855=>X"1B",
13856=>X"1B",
13857=>X"1B",
13858=>X"1B",
13859=>X"1A",
13860=>X"2A",
13861=>X"2F",
13862=>X"3E",
13863=>X"3E",
13864=>X"3A",
13865=>X"39",
13866=>X"38",
13867=>X"38",
13868=>X"38",
13869=>X"38",
13870=>X"38",
13871=>X"38",
13872=>X"38",
13873=>X"38",
13874=>X"38",
13875=>X"38",
13876=>X"38",
13877=>X"38",
13878=>X"38",
13879=>X"38",
13880=>X"38",
13881=>X"38",
13882=>X"29",
13883=>X"29",
13884=>X"15",
13885=>X"15",
13886=>X"15",
13887=>X"15",
13888=>X"15",
13889=>X"15",
13890=>X"15",
13891=>X"15",
13892=>X"15",
13893=>X"15",
13894=>X"15",
13895=>X"15",
13896=>X"15",
13897=>X"15",
13898=>X"15",
13899=>X"15",
13900=>X"15",
13901=>X"15",
13902=>X"15",
13903=>X"19",
13904=>X"19",
13905=>X"19",
13906=>X"19",
13907=>X"15",
13908=>X"15",
13909=>X"19",
13910=>X"15",
13911=>X"15",
13912=>X"15",
13913=>X"15",
13914=>X"15",
13915=>X"15",
13916=>X"15",
13917=>X"15",
13918=>X"15",
13919=>X"15",
13920=>X"15",
13921=>X"15",
13922=>X"15",
13923=>X"15",
13924=>X"00",
13925=>X"00",
13926=>X"00",
13927=>X"00",
13928=>X"00",
13929=>X"00",
13930=>X"00",
13931=>X"00",
13932=>X"00",
13933=>X"00",
13934=>X"00",
13935=>X"00",
13936=>X"00",
13937=>X"00",
13938=>X"00",
13939=>X"00",
13940=>X"00",
13941=>X"00",
13942=>X"00",
13943=>X"00",
13944=>X"00",
13945=>X"00",
13946=>X"00",
13947=>X"00",
13948=>X"00",
13949=>X"00",
13950=>X"00",
13951=>X"00",
13952=>X"00",
13953=>X"00",
13954=>X"00",
13955=>X"00",
13956=>X"00",
13957=>X"00",
13958=>X"00",
13959=>X"00",
13960=>X"00",
13961=>X"00",
13962=>X"00",
13963=>X"00",
13964=>X"00",
13965=>X"00",
13966=>X"00",
13967=>X"00",
13968=>X"00",
13969=>X"00",
13970=>X"00",
13971=>X"00",
13972=>X"00",
13973=>X"00",
13974=>X"00",
13975=>X"00",
13976=>X"00",
13977=>X"00",
13978=>X"00",
13979=>X"00",
13980=>X"00",
13981=>X"00",
13982=>X"00",
13983=>X"00",
13984=>X"00",
13985=>X"00",
13986=>X"00",
13987=>X"00",
13988=>X"00",
13989=>X"00",
13990=>X"00",
13991=>X"00",
13992=>X"00",
13993=>X"00",
13994=>X"00",
13995=>X"00",
13996=>X"00",
13997=>X"00",
13998=>X"00",
13999=>X"00",
14000=>X"00",
14001=>X"00",
14002=>X"00",
14003=>X"00",
14004=>X"00",
14005=>X"00",
14006=>X"00",
14007=>X"00",
14008=>X"00",
14009=>X"00",
14010=>X"00",
14011=>X"00",
14012=>X"00",
14013=>X"00",
14014=>X"00",
14015=>X"00",
14016=>X"00",
14017=>X"00",
14018=>X"00",
14019=>X"00",
14020=>X"00",
14021=>X"00",
14022=>X"00",
14023=>X"00",
14024=>X"00",
14025=>X"00",
14026=>X"00",
14027=>X"00",
14028=>X"00",
14029=>X"00",
14030=>X"00",
14031=>X"00",
14032=>X"00",
14033=>X"00",
14034=>X"00",
14035=>X"00",
14036=>X"00",
14037=>X"00",
14038=>X"00",
14039=>X"00",
14040=>X"00",
14041=>X"00",
14042=>X"00",
14043=>X"00",
14044=>X"00",
14045=>X"00",
14046=>X"00",
14047=>X"00",
14048=>X"00",
14049=>X"00",
14050=>X"00",
14051=>X"00",
14052=>X"00",
14053=>X"00",
14054=>X"00",
14055=>X"00",
14056=>X"00",
14057=>X"00",
14058=>X"00",
14059=>X"00",
14060=>X"00",
14061=>X"00",
14062=>X"00",
14063=>X"00",
14064=>X"00",
14065=>X"00",
14066=>X"00",
14067=>X"00",
14068=>X"00",
14069=>X"00",
14070=>X"00",
14071=>X"00",
14072=>X"00",
14073=>X"00",
14074=>X"00",
14075=>X"00",
14076=>X"00",
14077=>X"00",
14078=>X"00",
14079=>X"00",
14080=>X"14",
14081=>X"15",
14082=>X"15",
14083=>X"15",
14084=>X"15",
14085=>X"15",
14086=>X"15",
14087=>X"15",
14088=>X"15",
14089=>X"15",
14090=>X"14",
14091=>X"14",
14092=>X"14",
14093=>X"14",
14094=>X"14",
14095=>X"14",
14096=>X"14",
14097=>X"14",
14098=>X"14",
14099=>X"15",
14100=>X"15",
14101=>X"15",
14102=>X"16",
14103=>X"1A",
14104=>X"1B",
14105=>X"17",
14106=>X"17",
14107=>X"16",
14108=>X"16",
14109=>X"1B",
14110=>X"16",
14111=>X"16",
14112=>X"16",
14113=>X"1B",
14114=>X"1A",
14115=>X"16",
14116=>X"2A",
14117=>X"3E",
14118=>X"3E",
14119=>X"3A",
14120=>X"2E",
14121=>X"3D",
14122=>X"39",
14123=>X"3D",
14124=>X"38",
14125=>X"38",
14126=>X"38",
14127=>X"38",
14128=>X"38",
14129=>X"38",
14130=>X"38",
14131=>X"38",
14132=>X"38",
14133=>X"38",
14134=>X"38",
14135=>X"38",
14136=>X"28",
14137=>X"29",
14138=>X"25",
14139=>X"15",
14140=>X"15",
14141=>X"15",
14142=>X"15",
14143=>X"15",
14144=>X"15",
14145=>X"15",
14146=>X"15",
14147=>X"15",
14148=>X"15",
14149=>X"15",
14150=>X"15",
14151=>X"15",
14152=>X"15",
14153=>X"15",
14154=>X"15",
14155=>X"15",
14156=>X"15",
14157=>X"15",
14158=>X"15",
14159=>X"19",
14160=>X"19",
14161=>X"19",
14162=>X"15",
14163=>X"15",
14164=>X"15",
14165=>X"15",
14166=>X"15",
14167=>X"15",
14168=>X"15",
14169=>X"15",
14170=>X"15",
14171=>X"15",
14172=>X"15",
14173=>X"15",
14174=>X"15",
14175=>X"15",
14176=>X"15",
14177=>X"15",
14178=>X"15",
14179=>X"15",
14180=>X"00",
14181=>X"00",
14182=>X"00",
14183=>X"00",
14184=>X"00",
14185=>X"00",
14186=>X"00",
14187=>X"00",
14188=>X"00",
14189=>X"00",
14190=>X"00",
14191=>X"00",
14192=>X"00",
14193=>X"00",
14194=>X"00",
14195=>X"00",
14196=>X"00",
14197=>X"00",
14198=>X"00",
14199=>X"00",
14200=>X"00",
14201=>X"00",
14202=>X"00",
14203=>X"00",
14204=>X"00",
14205=>X"00",
14206=>X"00",
14207=>X"00",
14208=>X"00",
14209=>X"00",
14210=>X"00",
14211=>X"00",
14212=>X"00",
14213=>X"00",
14214=>X"00",
14215=>X"00",
14216=>X"00",
14217=>X"00",
14218=>X"00",
14219=>X"00",
14220=>X"00",
14221=>X"00",
14222=>X"00",
14223=>X"00",
14224=>X"00",
14225=>X"00",
14226=>X"00",
14227=>X"00",
14228=>X"00",
14229=>X"00",
14230=>X"00",
14231=>X"00",
14232=>X"00",
14233=>X"00",
14234=>X"00",
14235=>X"00",
14236=>X"00",
14237=>X"00",
14238=>X"00",
14239=>X"00",
14240=>X"00",
14241=>X"00",
14242=>X"00",
14243=>X"00",
14244=>X"00",
14245=>X"00",
14246=>X"00",
14247=>X"00",
14248=>X"00",
14249=>X"00",
14250=>X"00",
14251=>X"00",
14252=>X"00",
14253=>X"00",
14254=>X"00",
14255=>X"00",
14256=>X"00",
14257=>X"00",
14258=>X"00",
14259=>X"00",
14260=>X"00",
14261=>X"00",
14262=>X"00",
14263=>X"00",
14264=>X"00",
14265=>X"00",
14266=>X"00",
14267=>X"00",
14268=>X"00",
14269=>X"00",
14270=>X"00",
14271=>X"00",
14272=>X"00",
14273=>X"00",
14274=>X"00",
14275=>X"00",
14276=>X"00",
14277=>X"00",
14278=>X"00",
14279=>X"00",
14280=>X"00",
14281=>X"00",
14282=>X"00",
14283=>X"00",
14284=>X"00",
14285=>X"00",
14286=>X"00",
14287=>X"00",
14288=>X"00",
14289=>X"00",
14290=>X"00",
14291=>X"00",
14292=>X"00",
14293=>X"00",
14294=>X"00",
14295=>X"00",
14296=>X"00",
14297=>X"00",
14298=>X"00",
14299=>X"00",
14300=>X"00",
14301=>X"00",
14302=>X"00",
14303=>X"00",
14304=>X"00",
14305=>X"00",
14306=>X"00",
14307=>X"00",
14308=>X"00",
14309=>X"00",
14310=>X"00",
14311=>X"00",
14312=>X"00",
14313=>X"00",
14314=>X"00",
14315=>X"00",
14316=>X"00",
14317=>X"00",
14318=>X"00",
14319=>X"00",
14320=>X"00",
14321=>X"00",
14322=>X"00",
14323=>X"00",
14324=>X"00",
14325=>X"00",
14326=>X"00",
14327=>X"00",
14328=>X"00",
14329=>X"00",
14330=>X"00",
14331=>X"00",
14332=>X"00",
14333=>X"00",
14334=>X"00",
14335=>X"00",
14336=>X"04",
14337=>X"04",
14338=>X"15",
14339=>X"15",
14340=>X"15",
14341=>X"15",
14342=>X"15",
14343=>X"15",
14344=>X"15",
14345=>X"15",
14346=>X"14",
14347=>X"14",
14348=>X"14",
14349=>X"14",
14350=>X"14",
14351=>X"14",
14352=>X"14",
14353=>X"14",
14354=>X"15",
14355=>X"15",
14356=>X"16",
14357=>X"16",
14358=>X"16",
14359=>X"1B",
14360=>X"16",
14361=>X"17",
14362=>X"1A",
14363=>X"16",
14364=>X"16",
14365=>X"16",
14366=>X"16",
14367=>X"16",
14368=>X"16",
14369=>X"2A",
14370=>X"2A",
14371=>X"16",
14372=>X"2A",
14373=>X"2A",
14374=>X"3A",
14375=>X"2A",
14376=>X"3D",
14377=>X"39",
14378=>X"39",
14379=>X"29",
14380=>X"38",
14381=>X"28",
14382=>X"38",
14383=>X"28",
14384=>X"38",
14385=>X"38",
14386=>X"28",
14387=>X"38",
14388=>X"38",
14389=>X"28",
14390=>X"38",
14391=>X"28",
14392=>X"29",
14393=>X"25",
14394=>X"15",
14395=>X"15",
14396=>X"15",
14397=>X"15",
14398=>X"15",
14399=>X"15",
14400=>X"15",
14401=>X"15",
14402=>X"15",
14403=>X"15",
14404=>X"15",
14405=>X"15",
14406=>X"15",
14407=>X"15",
14408=>X"15",
14409=>X"15",
14410=>X"15",
14411=>X"15",
14412=>X"15",
14413=>X"19",
14414=>X"19",
14415=>X"15",
14416=>X"19",
14417=>X"25",
14418=>X"15",
14419=>X"19",
14420=>X"15",
14421=>X"15",
14422=>X"15",
14423=>X"15",
14424=>X"15",
14425=>X"15",
14426=>X"15",
14427=>X"15",
14428=>X"15",
14429=>X"15",
14430=>X"15",
14431=>X"15",
14432=>X"15",
14433=>X"15",
14434=>X"15",
14435=>X"15",
14436=>X"00",
14437=>X"00",
14438=>X"00",
14439=>X"00",
14440=>X"00",
14441=>X"00",
14442=>X"00",
14443=>X"00",
14444=>X"00",
14445=>X"00",
14446=>X"00",
14447=>X"00",
14448=>X"00",
14449=>X"00",
14450=>X"00",
14451=>X"00",
14452=>X"00",
14453=>X"00",
14454=>X"00",
14455=>X"00",
14456=>X"00",
14457=>X"00",
14458=>X"00",
14459=>X"00",
14460=>X"00",
14461=>X"00",
14462=>X"00",
14463=>X"00",
14464=>X"00",
14465=>X"00",
14466=>X"00",
14467=>X"00",
14468=>X"00",
14469=>X"00",
14470=>X"00",
14471=>X"00",
14472=>X"00",
14473=>X"00",
14474=>X"00",
14475=>X"00",
14476=>X"00",
14477=>X"00",
14478=>X"00",
14479=>X"00",
14480=>X"00",
14481=>X"00",
14482=>X"00",
14483=>X"00",
14484=>X"00",
14485=>X"00",
14486=>X"00",
14487=>X"00",
14488=>X"00",
14489=>X"00",
14490=>X"00",
14491=>X"00",
14492=>X"00",
14493=>X"00",
14494=>X"00",
14495=>X"00",
14496=>X"00",
14497=>X"00",
14498=>X"00",
14499=>X"00",
14500=>X"00",
14501=>X"00",
14502=>X"00",
14503=>X"00",
14504=>X"00",
14505=>X"00",
14506=>X"00",
14507=>X"00",
14508=>X"00",
14509=>X"00",
14510=>X"00",
14511=>X"00",
14512=>X"00",
14513=>X"00",
14514=>X"00",
14515=>X"00",
14516=>X"00",
14517=>X"00",
14518=>X"00",
14519=>X"00",
14520=>X"00",
14521=>X"00",
14522=>X"00",
14523=>X"00",
14524=>X"00",
14525=>X"00",
14526=>X"00",
14527=>X"00",
14528=>X"00",
14529=>X"00",
14530=>X"00",
14531=>X"00",
14532=>X"00",
14533=>X"00",
14534=>X"00",
14535=>X"00",
14536=>X"00",
14537=>X"00",
14538=>X"00",
14539=>X"00",
14540=>X"00",
14541=>X"00",
14542=>X"00",
14543=>X"00",
14544=>X"00",
14545=>X"00",
14546=>X"00",
14547=>X"00",
14548=>X"00",
14549=>X"00",
14550=>X"00",
14551=>X"00",
14552=>X"00",
14553=>X"00",
14554=>X"00",
14555=>X"00",
14556=>X"00",
14557=>X"00",
14558=>X"00",
14559=>X"00",
14560=>X"00",
14561=>X"00",
14562=>X"00",
14563=>X"00",
14564=>X"00",
14565=>X"00",
14566=>X"00",
14567=>X"00",
14568=>X"00",
14569=>X"00",
14570=>X"00",
14571=>X"00",
14572=>X"00",
14573=>X"00",
14574=>X"00",
14575=>X"00",
14576=>X"00",
14577=>X"00",
14578=>X"00",
14579=>X"00",
14580=>X"00",
14581=>X"00",
14582=>X"00",
14583=>X"00",
14584=>X"00",
14585=>X"00",
14586=>X"00",
14587=>X"00",
14588=>X"00",
14589=>X"00",
14590=>X"00",
14591=>X"00",
14592=>X"04",
14593=>X"04",
14594=>X"15",
14595=>X"15",
14596=>X"15",
14597=>X"15",
14598=>X"15",
14599=>X"15",
14600=>X"14",
14601=>X"14",
14602=>X"14",
14603=>X"14",
14604=>X"14",
14605=>X"14",
14606=>X"14",
14607=>X"14",
14608=>X"14",
14609=>X"14",
14610=>X"15",
14611=>X"15",
14612=>X"16",
14613=>X"16",
14614=>X"16",
14615=>X"16",
14616=>X"16",
14617=>X"16",
14618=>X"16",
14619=>X"16",
14620=>X"15",
14621=>X"15",
14622=>X"15",
14623=>X"15",
14624=>X"2A",
14625=>X"2A",
14626=>X"25",
14627=>X"25",
14628=>X"2A",
14629=>X"2A",
14630=>X"2A",
14631=>X"2A",
14632=>X"39",
14633=>X"39",
14634=>X"39",
14635=>X"29",
14636=>X"38",
14637=>X"28",
14638=>X"28",
14639=>X"28",
14640=>X"28",
14641=>X"38",
14642=>X"28",
14643=>X"28",
14644=>X"38",
14645=>X"28",
14646=>X"28",
14647=>X"28",
14648=>X"29",
14649=>X"29",
14650=>X"15",
14651=>X"15",
14652=>X"15",
14653=>X"15",
14654=>X"15",
14655=>X"15",
14656=>X"15",
14657=>X"15",
14658=>X"15",
14659=>X"15",
14660=>X"15",
14661=>X"15",
14662=>X"15",
14663=>X"15",
14664=>X"15",
14665=>X"15",
14666=>X"15",
14667=>X"15",
14668=>X"15",
14669=>X"15",
14670=>X"19",
14671=>X"19",
14672=>X"15",
14673=>X"15",
14674=>X"15",
14675=>X"15",
14676=>X"15",
14677=>X"15",
14678=>X"15",
14679=>X"15",
14680=>X"15",
14681=>X"15",
14682=>X"15",
14683=>X"15",
14684=>X"15",
14685=>X"15",
14686=>X"15",
14687=>X"15",
14688=>X"15",
14689=>X"15",
14690=>X"15",
14691=>X"15",
14692=>X"00",
14693=>X"00",
14694=>X"00",
14695=>X"00",
14696=>X"00",
14697=>X"00",
14698=>X"00",
14699=>X"00",
14700=>X"00",
14701=>X"00",
14702=>X"00",
14703=>X"00",
14704=>X"00",
14705=>X"00",
14706=>X"00",
14707=>X"00",
14708=>X"00",
14709=>X"00",
14710=>X"00",
14711=>X"00",
14712=>X"00",
14713=>X"00",
14714=>X"00",
14715=>X"00",
14716=>X"00",
14717=>X"00",
14718=>X"00",
14719=>X"00",
14720=>X"00",
14721=>X"00",
14722=>X"00",
14723=>X"00",
14724=>X"00",
14725=>X"00",
14726=>X"00",
14727=>X"00",
14728=>X"00",
14729=>X"00",
14730=>X"00",
14731=>X"00",
14732=>X"00",
14733=>X"00",
14734=>X"00",
14735=>X"00",
14736=>X"00",
14737=>X"00",
14738=>X"00",
14739=>X"00",
14740=>X"00",
14741=>X"00",
14742=>X"00",
14743=>X"00",
14744=>X"00",
14745=>X"00",
14746=>X"00",
14747=>X"00",
14748=>X"00",
14749=>X"00",
14750=>X"00",
14751=>X"00",
14752=>X"00",
14753=>X"00",
14754=>X"00",
14755=>X"00",
14756=>X"00",
14757=>X"00",
14758=>X"00",
14759=>X"00",
14760=>X"00",
14761=>X"00",
14762=>X"00",
14763=>X"00",
14764=>X"00",
14765=>X"00",
14766=>X"00",
14767=>X"00",
14768=>X"00",
14769=>X"00",
14770=>X"00",
14771=>X"00",
14772=>X"00",
14773=>X"00",
14774=>X"00",
14775=>X"00",
14776=>X"00",
14777=>X"00",
14778=>X"00",
14779=>X"00",
14780=>X"00",
14781=>X"00",
14782=>X"00",
14783=>X"00",
14784=>X"00",
14785=>X"00",
14786=>X"00",
14787=>X"00",
14788=>X"00",
14789=>X"00",
14790=>X"00",
14791=>X"00",
14792=>X"00",
14793=>X"00",
14794=>X"00",
14795=>X"00",
14796=>X"00",
14797=>X"00",
14798=>X"00",
14799=>X"00",
14800=>X"00",
14801=>X"00",
14802=>X"00",
14803=>X"00",
14804=>X"00",
14805=>X"00",
14806=>X"00",
14807=>X"00",
14808=>X"00",
14809=>X"00",
14810=>X"00",
14811=>X"00",
14812=>X"00",
14813=>X"00",
14814=>X"00",
14815=>X"00",
14816=>X"00",
14817=>X"00",
14818=>X"00",
14819=>X"00",
14820=>X"00",
14821=>X"00",
14822=>X"00",
14823=>X"00",
14824=>X"00",
14825=>X"00",
14826=>X"00",
14827=>X"00",
14828=>X"00",
14829=>X"00",
14830=>X"00",
14831=>X"00",
14832=>X"00",
14833=>X"00",
14834=>X"00",
14835=>X"00",
14836=>X"00",
14837=>X"00",
14838=>X"00",
14839=>X"00",
14840=>X"00",
14841=>X"00",
14842=>X"00",
14843=>X"00",
14844=>X"00",
14845=>X"00",
14846=>X"00",
14847=>X"00",
14848=>X"04",
14849=>X"04",
14850=>X"04",
14851=>X"04",
14852=>X"04",
14853=>X"05",
14854=>X"15",
14855=>X"15",
14856=>X"14",
14857=>X"14",
14858=>X"14",
14859=>X"14",
14860=>X"14",
14861=>X"14",
14862=>X"14",
14863=>X"14",
14864=>X"14",
14865=>X"15",
14866=>X"15",
14867=>X"15",
14868=>X"1A",
14869=>X"1B",
14870=>X"16",
14871=>X"16",
14872=>X"16",
14873=>X"16",
14874=>X"16",
14875=>X"16",
14876=>X"15",
14877=>X"15",
14878=>X"15",
14879=>X"25",
14880=>X"29",
14881=>X"15",
14882=>X"15",
14883=>X"25",
14884=>X"29",
14885=>X"29",
14886=>X"29",
14887=>X"29",
14888=>X"29",
14889=>X"29",
14890=>X"29",
14891=>X"29",
14892=>X"29",
14893=>X"28",
14894=>X"28",
14895=>X"24",
14896=>X"28",
14897=>X"24",
14898=>X"28",
14899=>X"28",
14900=>X"28",
14901=>X"28",
14902=>X"29",
14903=>X"15",
14904=>X"15",
14905=>X"15",
14906=>X"15",
14907=>X"15",
14908=>X"15",
14909=>X"15",
14910=>X"15",
14911=>X"15",
14912=>X"15",
14913=>X"15",
14914=>X"15",
14915=>X"15",
14916=>X"15",
14917=>X"15",
14918=>X"15",
14919=>X"15",
14920=>X"19",
14921=>X"19",
14922=>X"15",
14923=>X"15",
14924=>X"19",
14925=>X"15",
14926=>X"15",
14927=>X"15",
14928=>X"15",
14929=>X"15",
14930=>X"15",
14931=>X"15",
14932=>X"15",
14933=>X"15",
14934=>X"15",
14935=>X"15",
14936=>X"15",
14937=>X"15",
14938=>X"15",
14939=>X"15",
14940=>X"15",
14941=>X"15",
14942=>X"15",
14943=>X"15",
14944=>X"15",
14945=>X"15",
14946=>X"15",
14947=>X"15",
14948=>X"00",
14949=>X"00",
14950=>X"00",
14951=>X"00",
14952=>X"00",
14953=>X"00",
14954=>X"00",
14955=>X"00",
14956=>X"00",
14957=>X"00",
14958=>X"00",
14959=>X"00",
14960=>X"00",
14961=>X"00",
14962=>X"00",
14963=>X"00",
14964=>X"00",
14965=>X"00",
14966=>X"00",
14967=>X"00",
14968=>X"00",
14969=>X"00",
14970=>X"00",
14971=>X"00",
14972=>X"00",
14973=>X"00",
14974=>X"00",
14975=>X"00",
14976=>X"00",
14977=>X"00",
14978=>X"00",
14979=>X"00",
14980=>X"00",
14981=>X"00",
14982=>X"00",
14983=>X"00",
14984=>X"00",
14985=>X"00",
14986=>X"00",
14987=>X"00",
14988=>X"00",
14989=>X"00",
14990=>X"00",
14991=>X"00",
14992=>X"00",
14993=>X"00",
14994=>X"00",
14995=>X"00",
14996=>X"00",
14997=>X"00",
14998=>X"00",
14999=>X"00",
15000=>X"00",
15001=>X"00",
15002=>X"00",
15003=>X"00",
15004=>X"00",
15005=>X"00",
15006=>X"00",
15007=>X"00",
15008=>X"00",
15009=>X"00",
15010=>X"00",
15011=>X"00",
15012=>X"00",
15013=>X"00",
15014=>X"00",
15015=>X"00",
15016=>X"00",
15017=>X"00",
15018=>X"00",
15019=>X"00",
15020=>X"00",
15021=>X"00",
15022=>X"00",
15023=>X"00",
15024=>X"00",
15025=>X"00",
15026=>X"00",
15027=>X"00",
15028=>X"00",
15029=>X"00",
15030=>X"00",
15031=>X"00",
15032=>X"00",
15033=>X"00",
15034=>X"00",
15035=>X"00",
15036=>X"00",
15037=>X"00",
15038=>X"00",
15039=>X"00",
15040=>X"00",
15041=>X"00",
15042=>X"00",
15043=>X"00",
15044=>X"00",
15045=>X"00",
15046=>X"00",
15047=>X"00",
15048=>X"00",
15049=>X"00",
15050=>X"00",
15051=>X"00",
15052=>X"00",
15053=>X"00",
15054=>X"00",
15055=>X"00",
15056=>X"00",
15057=>X"00",
15058=>X"00",
15059=>X"00",
15060=>X"00",
15061=>X"00",
15062=>X"00",
15063=>X"00",
15064=>X"00",
15065=>X"00",
15066=>X"00",
15067=>X"00",
15068=>X"00",
15069=>X"00",
15070=>X"00",
15071=>X"00",
15072=>X"00",
15073=>X"00",
15074=>X"00",
15075=>X"00",
15076=>X"00",
15077=>X"00",
15078=>X"00",
15079=>X"00",
15080=>X"00",
15081=>X"00",
15082=>X"00",
15083=>X"00",
15084=>X"00",
15085=>X"00",
15086=>X"00",
15087=>X"00",
15088=>X"00",
15089=>X"00",
15090=>X"00",
15091=>X"00",
15092=>X"00",
15093=>X"00",
15094=>X"00",
15095=>X"00",
15096=>X"00",
15097=>X"00",
15098=>X"00",
15099=>X"00",
15100=>X"00",
15101=>X"00",
15102=>X"00",
15103=>X"00",
15104=>X"04",
15105=>X"04",
15106=>X"04",
15107=>X"14",
15108=>X"14",
15109=>X"14",
15110=>X"14",
15111=>X"14",
15112=>X"14",
15113=>X"14",
15114=>X"14",
15115=>X"14",
15116=>X"14",
15117=>X"14",
15118=>X"14",
15119=>X"14",
15120=>X"15",
15121=>X"15",
15122=>X"15",
15123=>X"16",
15124=>X"1B",
15125=>X"1B",
15126=>X"16",
15127=>X"16",
15128=>X"16",
15129=>X"16",
15130=>X"16",
15131=>X"16",
15132=>X"15",
15133=>X"15",
15134=>X"15",
15135=>X"15",
15136=>X"15",
15137=>X"15",
15138=>X"15",
15139=>X"15",
15140=>X"29",
15141=>X"29",
15142=>X"29",
15143=>X"29",
15144=>X"29",
15145=>X"29",
15146=>X"25",
15147=>X"25",
15148=>X"25",
15149=>X"25",
15150=>X"25",
15151=>X"24",
15152=>X"25",
15153=>X"25",
15154=>X"28",
15155=>X"28",
15156=>X"25",
15157=>X"25",
15158=>X"15",
15159=>X"15",
15160=>X"15",
15161=>X"15",
15162=>X"15",
15163=>X"15",
15164=>X"15",
15165=>X"15",
15166=>X"15",
15167=>X"15",
15168=>X"15",
15169=>X"15",
15170=>X"15",
15171=>X"15",
15172=>X"15",
15173=>X"15",
15174=>X"15",
15175=>X"15",
15176=>X"19",
15177=>X"19",
15178=>X"15",
15179=>X"15",
15180=>X"15",
15181=>X"15",
15182=>X"15",
15183=>X"15",
15184=>X"15",
15185=>X"15",
15186=>X"15",
15187=>X"15",
15188=>X"15",
15189=>X"15",
15190=>X"15",
15191=>X"15",
15192=>X"15",
15193=>X"15",
15194=>X"15",
15195=>X"15",
15196=>X"15",
15197=>X"15",
15198=>X"15",
15199=>X"15",
15200=>X"15",
15201=>X"15",
15202=>X"15",
15203=>X"15",
15204=>X"00",
15205=>X"00",
15206=>X"00",
15207=>X"00",
15208=>X"00",
15209=>X"00",
15210=>X"00",
15211=>X"00",
15212=>X"00",
15213=>X"00",
15214=>X"00",
15215=>X"00",
15216=>X"00",
15217=>X"00",
15218=>X"00",
15219=>X"00",
15220=>X"00",
15221=>X"00",
15222=>X"00",
15223=>X"00",
15224=>X"00",
15225=>X"00",
15226=>X"00",
15227=>X"00",
15228=>X"00",
15229=>X"00",
15230=>X"00",
15231=>X"00",
15232=>X"00",
15233=>X"00",
15234=>X"00",
15235=>X"00",
15236=>X"00",
15237=>X"00",
15238=>X"00",
15239=>X"00",
15240=>X"00",
15241=>X"00",
15242=>X"00",
15243=>X"00",
15244=>X"00",
15245=>X"00",
15246=>X"00",
15247=>X"00",
15248=>X"00",
15249=>X"00",
15250=>X"00",
15251=>X"00",
15252=>X"00",
15253=>X"00",
15254=>X"00",
15255=>X"00",
15256=>X"00",
15257=>X"00",
15258=>X"00",
15259=>X"00",
15260=>X"00",
15261=>X"00",
15262=>X"00",
15263=>X"00",
15264=>X"00",
15265=>X"00",
15266=>X"00",
15267=>X"00",
15268=>X"00",
15269=>X"00",
15270=>X"00",
15271=>X"00",
15272=>X"00",
15273=>X"00",
15274=>X"00",
15275=>X"00",
15276=>X"00",
15277=>X"00",
15278=>X"00",
15279=>X"00",
15280=>X"00",
15281=>X"00",
15282=>X"00",
15283=>X"00",
15284=>X"00",
15285=>X"00",
15286=>X"00",
15287=>X"00",
15288=>X"00",
15289=>X"00",
15290=>X"00",
15291=>X"00",
15292=>X"00",
15293=>X"00",
15294=>X"00",
15295=>X"00",
15296=>X"00",
15297=>X"00",
15298=>X"00",
15299=>X"00",
15300=>X"00",
15301=>X"00",
15302=>X"00",
15303=>X"00",
15304=>X"00",
15305=>X"00",
15306=>X"00",
15307=>X"00",
15308=>X"00",
15309=>X"00",
15310=>X"00",
15311=>X"00",
15312=>X"00",
15313=>X"00",
15314=>X"00",
15315=>X"00",
15316=>X"00",
15317=>X"00",
15318=>X"00",
15319=>X"00",
15320=>X"00",
15321=>X"00",
15322=>X"00",
15323=>X"00",
15324=>X"00",
15325=>X"00",
15326=>X"00",
15327=>X"00",
15328=>X"00",
15329=>X"00",
15330=>X"00",
15331=>X"00",
15332=>X"00",
15333=>X"00",
15334=>X"00",
15335=>X"00",
15336=>X"00",
15337=>X"00",
15338=>X"00",
15339=>X"00",
15340=>X"00",
15341=>X"00",
15342=>X"00",
15343=>X"00",
15344=>X"00",
15345=>X"00",
15346=>X"00",
15347=>X"00",
15348=>X"00",
15349=>X"00",
15350=>X"00",
15351=>X"00",
15352=>X"00",
15353=>X"00",
15354=>X"00",
15355=>X"00",
15356=>X"00",
15357=>X"00",
15358=>X"00",
15359=>X"00",
15360=>X"04",
15361=>X"04",
15362=>X"04",
15363=>X"14",
15364=>X"14",
15365=>X"14",
15366=>X"04",
15367=>X"14",
15368=>X"14",
15369=>X"14",
15370=>X"14",
15371=>X"14",
15372=>X"14",
15373=>X"14",
15374=>X"14",
15375=>X"14",
15376=>X"15",
15377=>X"15",
15378=>X"15",
15379=>X"16",
15380=>X"16",
15381=>X"16",
15382=>X"16",
15383=>X"16",
15384=>X"16",
15385=>X"16",
15386=>X"15",
15387=>X"15",
15388=>X"15",
15389=>X"15",
15390=>X"15",
15391=>X"15",
15392=>X"15",
15393=>X"15",
15394=>X"15",
15395=>X"15",
15396=>X"25",
15397=>X"25",
15398=>X"15",
15399=>X"15",
15400=>X"15",
15401=>X"15",
15402=>X"15",
15403=>X"15",
15404=>X"15",
15405=>X"25",
15406=>X"25",
15407=>X"25",
15408=>X"25",
15409=>X"25",
15410=>X"29",
15411=>X"25",
15412=>X"25",
15413=>X"15",
15414=>X"15",
15415=>X"15",
15416=>X"15",
15417=>X"15",
15418=>X"15",
15419=>X"15",
15420=>X"15",
15421=>X"15",
15422=>X"15",
15423=>X"15",
15424=>X"15",
15425=>X"15",
15426=>X"15",
15427=>X"15",
15428=>X"15",
15429=>X"15",
15430=>X"15",
15431=>X"15",
15432=>X"15",
15433=>X"15",
15434=>X"19",
15435=>X"15",
15436=>X"15",
15437=>X"15",
15438=>X"15",
15439=>X"15",
15440=>X"15",
15441=>X"15",
15442=>X"15",
15443=>X"15",
15444=>X"15",
15445=>X"15",
15446=>X"15",
15447=>X"15",
15448=>X"15",
15449=>X"15",
15450=>X"15",
15451=>X"15",
15452=>X"15",
15453=>X"15",
15454=>X"15",
15455=>X"15",
15456=>X"15",
15457=>X"15",
15458=>X"15",
15459=>X"15",
15460=>X"00",
15461=>X"00",
15462=>X"00",
15463=>X"00",
15464=>X"00",
15465=>X"00",
15466=>X"00",
15467=>X"00",
15468=>X"00",
15469=>X"00",
15470=>X"00",
15471=>X"00",
15472=>X"00",
15473=>X"00",
15474=>X"00",
15475=>X"00",
15476=>X"00",
15477=>X"00",
15478=>X"00",
15479=>X"00",
15480=>X"00",
15481=>X"00",
15482=>X"00",
15483=>X"00",
15484=>X"00",
15485=>X"00",
15486=>X"00",
15487=>X"00",
15488=>X"00",
15489=>X"00",
15490=>X"00",
15491=>X"00",
15492=>X"00",
15493=>X"00",
15494=>X"00",
15495=>X"00",
15496=>X"00",
15497=>X"00",
15498=>X"00",
15499=>X"00",
15500=>X"00",
15501=>X"00",
15502=>X"00",
15503=>X"00",
15504=>X"00",
15505=>X"00",
15506=>X"00",
15507=>X"00",
15508=>X"00",
15509=>X"00",
15510=>X"00",
15511=>X"00",
15512=>X"00",
15513=>X"00",
15514=>X"00",
15515=>X"00",
15516=>X"00",
15517=>X"00",
15518=>X"00",
15519=>X"00",
15520=>X"00",
15521=>X"00",
15522=>X"00",
15523=>X"00",
15524=>X"00",
15525=>X"00",
15526=>X"00",
15527=>X"00",
15528=>X"00",
15529=>X"00",
15530=>X"00",
15531=>X"00",
15532=>X"00",
15533=>X"00",
15534=>X"00",
15535=>X"00",
15536=>X"00",
15537=>X"00",
15538=>X"00",
15539=>X"00",
15540=>X"00",
15541=>X"00",
15542=>X"00",
15543=>X"00",
15544=>X"00",
15545=>X"00",
15546=>X"00",
15547=>X"00",
15548=>X"00",
15549=>X"00",
15550=>X"00",
15551=>X"00",
15552=>X"00",
15553=>X"00",
15554=>X"00",
15555=>X"00",
15556=>X"00",
15557=>X"00",
15558=>X"00",
15559=>X"00",
15560=>X"00",
15561=>X"00",
15562=>X"00",
15563=>X"00",
15564=>X"00",
15565=>X"00",
15566=>X"00",
15567=>X"00",
15568=>X"00",
15569=>X"00",
15570=>X"00",
15571=>X"00",
15572=>X"00",
15573=>X"00",
15574=>X"00",
15575=>X"00",
15576=>X"00",
15577=>X"00",
15578=>X"00",
15579=>X"00",
15580=>X"00",
15581=>X"00",
15582=>X"00",
15583=>X"00",
15584=>X"00",
15585=>X"00",
15586=>X"00",
15587=>X"00",
15588=>X"00",
15589=>X"00",
15590=>X"00",
15591=>X"00",
15592=>X"00",
15593=>X"00",
15594=>X"00",
15595=>X"00",
15596=>X"00",
15597=>X"00",
15598=>X"00",
15599=>X"00",
15600=>X"00",
15601=>X"00",
15602=>X"00",
15603=>X"00",
15604=>X"00",
15605=>X"00",
15606=>X"00",
15607=>X"00",
15608=>X"00",
15609=>X"00",
15610=>X"00",
15611=>X"00",
15612=>X"00",
15613=>X"00",
15614=>X"00",
15615=>X"00",
15616=>X"04",
15617=>X"04",
15618=>X"04",
15619=>X"14",
15620=>X"14",
15621=>X"14",
15622=>X"04",
15623=>X"14",
15624=>X"14",
15625=>X"14",
15626=>X"14",
15627=>X"14",
15628=>X"14",
15629=>X"14",
15630=>X"14",
15631=>X"14",
15632=>X"15",
15633=>X"15",
15634=>X"15",
15635=>X"16",
15636=>X"16",
15637=>X"16",
15638=>X"16",
15639=>X"16",
15640=>X"16",
15641=>X"16",
15642=>X"15",
15643=>X"15",
15644=>X"15",
15645=>X"25",
15646=>X"15",
15647=>X"15",
15648=>X"15",
15649=>X"15",
15650=>X"15",
15651=>X"15",
15652=>X"25",
15653=>X"25",
15654=>X"15",
15655=>X"15",
15656=>X"25",
15657=>X"15",
15658=>X"15",
15659=>X"15",
15660=>X"15",
15661=>X"25",
15662=>X"25",
15663=>X"25",
15664=>X"15",
15665=>X"29",
15666=>X"25",
15667=>X"25",
15668=>X"15",
15669=>X"15",
15670=>X"15",
15671=>X"15",
15672=>X"15",
15673=>X"15",
15674=>X"15",
15675=>X"15",
15676=>X"15",
15677=>X"15",
15678=>X"15",
15679=>X"15",
15680=>X"15",
15681=>X"15",
15682=>X"15",
15683=>X"15",
15684=>X"15",
15685=>X"15",
15686=>X"15",
15687=>X"15",
15688=>X"15",
15689=>X"15",
15690=>X"15",
15691=>X"15",
15692=>X"15",
15693=>X"15",
15694=>X"15",
15695=>X"15",
15696=>X"15",
15697=>X"15",
15698=>X"15",
15699=>X"15",
15700=>X"15",
15701=>X"15",
15702=>X"15",
15703=>X"15",
15704=>X"15",
15705=>X"15",
15706=>X"15",
15707=>X"15",
15708=>X"15",
15709=>X"15",
15710=>X"15",
15711=>X"15",
15712=>X"15",
15713=>X"15",
15714=>X"15",
15715=>X"15",
15716=>X"00",
15717=>X"00",
15718=>X"00",
15719=>X"00",
15720=>X"00",
15721=>X"00",
15722=>X"00",
15723=>X"00",
15724=>X"00",
15725=>X"00",
15726=>X"00",
15727=>X"00",
15728=>X"00",
15729=>X"00",
15730=>X"00",
15731=>X"00",
15732=>X"00",
15733=>X"00",
15734=>X"00",
15735=>X"00",
15736=>X"00",
15737=>X"00",
15738=>X"00",
15739=>X"00",
15740=>X"00",
15741=>X"00",
15742=>X"00",
15743=>X"00",
15744=>X"00",
15745=>X"00",
15746=>X"00",
15747=>X"00",
15748=>X"00",
15749=>X"00",
15750=>X"00",
15751=>X"00",
15752=>X"00",
15753=>X"00",
15754=>X"00",
15755=>X"00",
15756=>X"00",
15757=>X"00",
15758=>X"00",
15759=>X"00",
15760=>X"00",
15761=>X"00",
15762=>X"00",
15763=>X"00",
15764=>X"00",
15765=>X"00",
15766=>X"00",
15767=>X"00",
15768=>X"00",
15769=>X"00",
15770=>X"00",
15771=>X"00",
15772=>X"00",
15773=>X"00",
15774=>X"00",
15775=>X"00",
15776=>X"00",
15777=>X"00",
15778=>X"00",
15779=>X"00",
15780=>X"00",
15781=>X"00",
15782=>X"00",
15783=>X"00",
15784=>X"00",
15785=>X"00",
15786=>X"00",
15787=>X"00",
15788=>X"00",
15789=>X"00",
15790=>X"00",
15791=>X"00",
15792=>X"00",
15793=>X"00",
15794=>X"00",
15795=>X"00",
15796=>X"00",
15797=>X"00",
15798=>X"00",
15799=>X"00",
15800=>X"00",
15801=>X"00",
15802=>X"00",
15803=>X"00",
15804=>X"00",
15805=>X"00",
15806=>X"00",
15807=>X"00",
15808=>X"00",
15809=>X"00",
15810=>X"00",
15811=>X"00",
15812=>X"00",
15813=>X"00",
15814=>X"00",
15815=>X"00",
15816=>X"00",
15817=>X"00",
15818=>X"00",
15819=>X"00",
15820=>X"00",
15821=>X"00",
15822=>X"00",
15823=>X"00",
15824=>X"00",
15825=>X"00",
15826=>X"00",
15827=>X"00",
15828=>X"00",
15829=>X"00",
15830=>X"00",
15831=>X"00",
15832=>X"00",
15833=>X"00",
15834=>X"00",
15835=>X"00",
15836=>X"00",
15837=>X"00",
15838=>X"00",
15839=>X"00",
15840=>X"00",
15841=>X"00",
15842=>X"00",
15843=>X"00",
15844=>X"00",
15845=>X"00",
15846=>X"00",
15847=>X"00",
15848=>X"00",
15849=>X"00",
15850=>X"00",
15851=>X"00",
15852=>X"00",
15853=>X"00",
15854=>X"00",
15855=>X"00",
15856=>X"00",
15857=>X"00",
15858=>X"00",
15859=>X"00",
15860=>X"00",
15861=>X"00",
15862=>X"00",
15863=>X"00",
15864=>X"00",
15865=>X"00",
15866=>X"00",
15867=>X"00",
15868=>X"00",
15869=>X"00",
15870=>X"00",
15871=>X"00",
15872=>X"04",
15873=>X"04",
15874=>X"04",
15875=>X"04",
15876=>X"05",
15877=>X"05",
15878=>X"04",
15879=>X"14",
15880=>X"14",
15881=>X"14",
15882=>X"04",
15883=>X"04",
15884=>X"14",
15885=>X"14",
15886=>X"14",
15887=>X"15",
15888=>X"15",
15889=>X"15",
15890=>X"15",
15891=>X"16",
15892=>X"17",
15893=>X"17",
15894=>X"16",
15895=>X"16",
15896=>X"16",
15897=>X"16",
15898=>X"15",
15899=>X"15",
15900=>X"25",
15901=>X"25",
15902=>X"15",
15903=>X"15",
15904=>X"15",
15905=>X"15",
15906=>X"15",
15907=>X"15",
15908=>X"15",
15909=>X"15",
15910=>X"15",
15911=>X"15",
15912=>X"15",
15913=>X"15",
15914=>X"15",
15915=>X"15",
15916=>X"25",
15917=>X"25",
15918=>X"25",
15919=>X"25",
15920=>X"15",
15921=>X"15",
15922=>X"15",
15923=>X"15",
15924=>X"15",
15925=>X"15",
15926=>X"15",
15927=>X"15",
15928=>X"15",
15929=>X"15",
15930=>X"15",
15931=>X"15",
15932=>X"15",
15933=>X"15",
15934=>X"15",
15935=>X"15",
15936=>X"15",
15937=>X"15",
15938=>X"15",
15939=>X"15",
15940=>X"15",
15941=>X"15",
15942=>X"15",
15943=>X"15",
15944=>X"15",
15945=>X"15",
15946=>X"15",
15947=>X"15",
15948=>X"15",
15949=>X"15",
15950=>X"15",
15951=>X"15",
15952=>X"15",
15953=>X"15",
15954=>X"15",
15955=>X"15",
15956=>X"15",
15957=>X"15",
15958=>X"15",
15959=>X"15",
15960=>X"15",
15961=>X"15",
15962=>X"15",
15963=>X"15",
15964=>X"15",
15965=>X"15",
15966=>X"15",
15967=>X"15",
15968=>X"15",
15969=>X"15",
15970=>X"15",
15971=>X"15",
15972=>X"00",
15973=>X"00",
15974=>X"00",
15975=>X"00",
15976=>X"00",
15977=>X"00",
15978=>X"00",
15979=>X"00",
15980=>X"00",
15981=>X"00",
15982=>X"00",
15983=>X"00",
15984=>X"00",
15985=>X"00",
15986=>X"00",
15987=>X"00",
15988=>X"00",
15989=>X"00",
15990=>X"00",
15991=>X"00",
15992=>X"00",
15993=>X"00",
15994=>X"00",
15995=>X"00",
15996=>X"00",
15997=>X"00",
15998=>X"00",
15999=>X"00",
16000=>X"00",
16001=>X"00",
16002=>X"00",
16003=>X"00",
16004=>X"00",
16005=>X"00",
16006=>X"00",
16007=>X"00",
16008=>X"00",
16009=>X"00",
16010=>X"00",
16011=>X"00",
16012=>X"00",
16013=>X"00",
16014=>X"00",
16015=>X"00",
16016=>X"00",
16017=>X"00",
16018=>X"00",
16019=>X"00",
16020=>X"00",
16021=>X"00",
16022=>X"00",
16023=>X"00",
16024=>X"00",
16025=>X"00",
16026=>X"00",
16027=>X"00",
16028=>X"00",
16029=>X"00",
16030=>X"00",
16031=>X"00",
16032=>X"00",
16033=>X"00",
16034=>X"00",
16035=>X"00",
16036=>X"00",
16037=>X"00",
16038=>X"00",
16039=>X"00",
16040=>X"00",
16041=>X"00",
16042=>X"00",
16043=>X"00",
16044=>X"00",
16045=>X"00",
16046=>X"00",
16047=>X"00",
16048=>X"00",
16049=>X"00",
16050=>X"00",
16051=>X"00",
16052=>X"00",
16053=>X"00",
16054=>X"00",
16055=>X"00",
16056=>X"00",
16057=>X"00",
16058=>X"00",
16059=>X"00",
16060=>X"00",
16061=>X"00",
16062=>X"00",
16063=>X"00",
16064=>X"00",
16065=>X"00",
16066=>X"00",
16067=>X"00",
16068=>X"00",
16069=>X"00",
16070=>X"00",
16071=>X"00",
16072=>X"00",
16073=>X"00",
16074=>X"00",
16075=>X"00",
16076=>X"00",
16077=>X"00",
16078=>X"00",
16079=>X"00",
16080=>X"00",
16081=>X"00",
16082=>X"00",
16083=>X"00",
16084=>X"00",
16085=>X"00",
16086=>X"00",
16087=>X"00",
16088=>X"00",
16089=>X"00",
16090=>X"00",
16091=>X"00",
16092=>X"00",
16093=>X"00",
16094=>X"00",
16095=>X"00",
16096=>X"00",
16097=>X"00",
16098=>X"00",
16099=>X"00",
16100=>X"00",
16101=>X"00",
16102=>X"00",
16103=>X"00",
16104=>X"00",
16105=>X"00",
16106=>X"00",
16107=>X"00",
16108=>X"00",
16109=>X"00",
16110=>X"00",
16111=>X"00",
16112=>X"00",
16113=>X"00",
16114=>X"00",
16115=>X"00",
16116=>X"00",
16117=>X"00",
16118=>X"00",
16119=>X"00",
16120=>X"00",
16121=>X"00",
16122=>X"00",
16123=>X"00",
16124=>X"00",
16125=>X"00",
16126=>X"00",
16127=>X"00",
16128=>X"04",
16129=>X"04",
16130=>X"04",
16131=>X"05",
16132=>X"05",
16133=>X"05",
16134=>X"05",
16135=>X"05",
16136=>X"05",
16137=>X"04",
16138=>X"04",
16139=>X"04",
16140=>X"14",
16141=>X"14",
16142=>X"15",
16143=>X"15",
16144=>X"15",
16145=>X"15",
16146=>X"15",
16147=>X"16",
16148=>X"1B",
16149=>X"17",
16150=>X"16",
16151=>X"16",
16152=>X"16",
16153=>X"15",
16154=>X"15",
16155=>X"15",
16156=>X"25",
16157=>X"25",
16158=>X"15",
16159=>X"15",
16160=>X"15",
16161=>X"15",
16162=>X"15",
16163=>X"15",
16164=>X"15",
16165=>X"15",
16166=>X"15",
16167=>X"15",
16168=>X"15",
16169=>X"15",
16170=>X"15",
16171=>X"15",
16172=>X"15",
16173=>X"25",
16174=>X"25",
16175=>X"25",
16176=>X"29",
16177=>X"15",
16178=>X"15",
16179=>X"15",
16180=>X"15",
16181=>X"15",
16182=>X"15",
16183=>X"15",
16184=>X"15",
16185=>X"15",
16186=>X"15",
16187=>X"15",
16188=>X"15",
16189=>X"15",
16190=>X"15",
16191=>X"15",
16192=>X"15",
16193=>X"15",
16194=>X"15",
16195=>X"15",
16196=>X"15",
16197=>X"15",
16198=>X"15",
16199=>X"15",
16200=>X"15",
16201=>X"15",
16202=>X"15",
16203=>X"15",
16204=>X"15",
16205=>X"15",
16206=>X"15",
16207=>X"15",
16208=>X"15",
16209=>X"15",
16210=>X"15",
16211=>X"15",
16212=>X"15",
16213=>X"15",
16214=>X"15",
16215=>X"15",
16216=>X"15",
16217=>X"15",
16218=>X"15",
16219=>X"15",
16220=>X"15",
16221=>X"15",
16222=>X"15",
16223=>X"15",
16224=>X"15",
16225=>X"15",
16226=>X"15",
16227=>X"15",
16228=>X"00",
16229=>X"00",
16230=>X"00",
16231=>X"00",
16232=>X"00",
16233=>X"00",
16234=>X"00",
16235=>X"00",
16236=>X"00",
16237=>X"00",
16238=>X"00",
16239=>X"00",
16240=>X"00",
16241=>X"00",
16242=>X"00",
16243=>X"00",
16244=>X"00",
16245=>X"00",
16246=>X"00",
16247=>X"00",
16248=>X"00",
16249=>X"00",
16250=>X"00",
16251=>X"00",
16252=>X"00",
16253=>X"00",
16254=>X"00",
16255=>X"00",
16256=>X"00",
16257=>X"00",
16258=>X"00",
16259=>X"00",
16260=>X"00",
16261=>X"00",
16262=>X"00",
16263=>X"00",
16264=>X"00",
16265=>X"00",
16266=>X"00",
16267=>X"00",
16268=>X"00",
16269=>X"00",
16270=>X"00",
16271=>X"00",
16272=>X"00",
16273=>X"00",
16274=>X"00",
16275=>X"00",
16276=>X"00",
16277=>X"00",
16278=>X"00",
16279=>X"00",
16280=>X"00",
16281=>X"00",
16282=>X"00",
16283=>X"00",
16284=>X"00",
16285=>X"00",
16286=>X"00",
16287=>X"00",
16288=>X"00",
16289=>X"00",
16290=>X"00",
16291=>X"00",
16292=>X"00",
16293=>X"00",
16294=>X"00",
16295=>X"00",
16296=>X"00",
16297=>X"00",
16298=>X"00",
16299=>X"00",
16300=>X"00",
16301=>X"00",
16302=>X"00",
16303=>X"00",
16304=>X"00",
16305=>X"00",
16306=>X"00",
16307=>X"00",
16308=>X"00",
16309=>X"00",
16310=>X"00",
16311=>X"00",
16312=>X"00",
16313=>X"00",
16314=>X"00",
16315=>X"00",
16316=>X"00",
16317=>X"00",
16318=>X"00",
16319=>X"00",
16320=>X"00",
16321=>X"00",
16322=>X"00",
16323=>X"00",
16324=>X"00",
16325=>X"00",
16326=>X"00",
16327=>X"00",
16328=>X"00",
16329=>X"00",
16330=>X"00",
16331=>X"00",
16332=>X"00",
16333=>X"00",
16334=>X"00",
16335=>X"00",
16336=>X"00",
16337=>X"00",
16338=>X"00",
16339=>X"00",
16340=>X"00",
16341=>X"00",
16342=>X"00",
16343=>X"00",
16344=>X"00",
16345=>X"00",
16346=>X"00",
16347=>X"00",
16348=>X"00",
16349=>X"00",
16350=>X"00",
16351=>X"00",
16352=>X"00",
16353=>X"00",
16354=>X"00",
16355=>X"00",
16356=>X"00",
16357=>X"00",
16358=>X"00",
16359=>X"00",
16360=>X"00",
16361=>X"00",
16362=>X"00",
16363=>X"00",
16364=>X"00",
16365=>X"00",
16366=>X"00",
16367=>X"00",
16368=>X"00",
16369=>X"00",
16370=>X"00",
16371=>X"00",
16372=>X"00",
16373=>X"00",
16374=>X"00",
16375=>X"00",
16376=>X"00",
16377=>X"00",
16378=>X"00",
16379=>X"00",
16380=>X"00",
16381=>X"00",
16382=>X"00",
16383=>X"00",
16384=>X"04",
16385=>X"04",
16386=>X"04",
16387=>X"05",
16388=>X"05",
16389=>X"05",
16390=>X"15",
16391=>X"15",
16392=>X"15",
16393=>X"04",
16394=>X"04",
16395=>X"04",
16396=>X"14",
16397=>X"15",
16398=>X"15",
16399=>X"15",
16400=>X"15",
16401=>X"15",
16402=>X"15",
16403=>X"16",
16404=>X"1A",
16405=>X"1A",
16406=>X"15",
16407=>X"15",
16408=>X"15",
16409=>X"15",
16410=>X"15",
16411=>X"15",
16412=>X"25",
16413=>X"25",
16414=>X"15",
16415=>X"15",
16416=>X"15",
16417=>X"15",
16418=>X"15",
16419=>X"15",
16420=>X"15",
16421=>X"15",
16422=>X"15",
16423=>X"15",
16424=>X"15",
16425=>X"15",
16426=>X"15",
16427=>X"15",
16428=>X"15",
16429=>X"15",
16430=>X"15",
16431=>X"25",
16432=>X"39",
16433=>X"2A",
16434=>X"25",
16435=>X"15",
16436=>X"15",
16437=>X"15",
16438=>X"15",
16439=>X"15",
16440=>X"15",
16441=>X"15",
16442=>X"15",
16443=>X"15",
16444=>X"15",
16445=>X"15",
16446=>X"15",
16447=>X"15",
16448=>X"15",
16449=>X"15",
16450=>X"15",
16451=>X"15",
16452=>X"15",
16453=>X"15",
16454=>X"15",
16455=>X"15",
16456=>X"15",
16457=>X"15",
16458=>X"15",
16459=>X"15",
16460=>X"15",
16461=>X"15",
16462=>X"15",
16463=>X"15",
16464=>X"15",
16465=>X"15",
16466=>X"15",
16467=>X"15",
16468=>X"15",
16469=>X"15",
16470=>X"15",
16471=>X"15",
16472=>X"15",
16473=>X"15",
16474=>X"15",
16475=>X"15",
16476=>X"15",
16477=>X"15",
16478=>X"15",
16479=>X"15",
16480=>X"15",
16481=>X"15",
16482=>X"15",
16483=>X"15",
16484=>X"00",
16485=>X"00",
16486=>X"00",
16487=>X"00",
16488=>X"00",
16489=>X"00",
16490=>X"00",
16491=>X"00",
16492=>X"00",
16493=>X"00",
16494=>X"00",
16495=>X"00",
16496=>X"00",
16497=>X"00",
16498=>X"00",
16499=>X"00",
16500=>X"00",
16501=>X"00",
16502=>X"00",
16503=>X"00",
16504=>X"00",
16505=>X"00",
16506=>X"00",
16507=>X"00",
16508=>X"00",
16509=>X"00",
16510=>X"00",
16511=>X"00",
16512=>X"00",
16513=>X"00",
16514=>X"00",
16515=>X"00",
16516=>X"00",
16517=>X"00",
16518=>X"00",
16519=>X"00",
16520=>X"00",
16521=>X"00",
16522=>X"00",
16523=>X"00",
16524=>X"00",
16525=>X"00",
16526=>X"00",
16527=>X"00",
16528=>X"00",
16529=>X"00",
16530=>X"00",
16531=>X"00",
16532=>X"00",
16533=>X"00",
16534=>X"00",
16535=>X"00",
16536=>X"00",
16537=>X"00",
16538=>X"00",
16539=>X"00",
16540=>X"00",
16541=>X"00",
16542=>X"00",
16543=>X"00",
16544=>X"00",
16545=>X"00",
16546=>X"00",
16547=>X"00",
16548=>X"00",
16549=>X"00",
16550=>X"00",
16551=>X"00",
16552=>X"00",
16553=>X"00",
16554=>X"00",
16555=>X"00",
16556=>X"00",
16557=>X"00",
16558=>X"00",
16559=>X"00",
16560=>X"00",
16561=>X"00",
16562=>X"00",
16563=>X"00",
16564=>X"00",
16565=>X"00",
16566=>X"00",
16567=>X"00",
16568=>X"00",
16569=>X"00",
16570=>X"00",
16571=>X"00",
16572=>X"00",
16573=>X"00",
16574=>X"00",
16575=>X"00",
16576=>X"00",
16577=>X"00",
16578=>X"00",
16579=>X"00",
16580=>X"00",
16581=>X"00",
16582=>X"00",
16583=>X"00",
16584=>X"00",
16585=>X"00",
16586=>X"00",
16587=>X"00",
16588=>X"00",
16589=>X"00",
16590=>X"00",
16591=>X"00",
16592=>X"00",
16593=>X"00",
16594=>X"00",
16595=>X"00",
16596=>X"00",
16597=>X"00",
16598=>X"00",
16599=>X"00",
16600=>X"00",
16601=>X"00",
16602=>X"00",
16603=>X"00",
16604=>X"00",
16605=>X"00",
16606=>X"00",
16607=>X"00",
16608=>X"00",
16609=>X"00",
16610=>X"00",
16611=>X"00",
16612=>X"00",
16613=>X"00",
16614=>X"00",
16615=>X"00",
16616=>X"00",
16617=>X"00",
16618=>X"00",
16619=>X"00",
16620=>X"00",
16621=>X"00",
16622=>X"00",
16623=>X"00",
16624=>X"00",
16625=>X"00",
16626=>X"00",
16627=>X"00",
16628=>X"00",
16629=>X"00",
16630=>X"00",
16631=>X"00",
16632=>X"00",
16633=>X"00",
16634=>X"00",
16635=>X"00",
16636=>X"00",
16637=>X"00",
16638=>X"00",
16639=>X"00",
16640=>X"04",
16641=>X"04",
16642=>X"04",
16643=>X"04",
16644=>X"04",
16645=>X"04",
16646=>X"14",
16647=>X"14",
16648=>X"14",
16649=>X"04",
16650=>X"04",
16651=>X"04",
16652=>X"15",
16653=>X"15",
16654=>X"15",
16655=>X"15",
16656=>X"15",
16657=>X"15",
16658=>X"15",
16659=>X"15",
16660=>X"1A",
16661=>X"15",
16662=>X"15",
16663=>X"15",
16664=>X"15",
16665=>X"15",
16666=>X"29",
16667=>X"25",
16668=>X"25",
16669=>X"25",
16670=>X"15",
16671=>X"15",
16672=>X"15",
16673=>X"15",
16674=>X"15",
16675=>X"15",
16676=>X"15",
16677=>X"15",
16678=>X"15",
16679=>X"15",
16680=>X"15",
16681=>X"15",
16682=>X"15",
16683=>X"15",
16684=>X"15",
16685=>X"15",
16686=>X"29",
16687=>X"29",
16688=>X"3A",
16689=>X"3A",
16690=>X"3A",
16691=>X"26",
16692=>X"25",
16693=>X"15",
16694=>X"15",
16695=>X"15",
16696=>X"15",
16697=>X"15",
16698=>X"15",
16699=>X"15",
16700=>X"15",
16701=>X"15",
16702=>X"15",
16703=>X"15",
16704=>X"15",
16705=>X"15",
16706=>X"15",
16707=>X"15",
16708=>X"15",
16709=>X"15",
16710=>X"15",
16711=>X"15",
16712=>X"15",
16713=>X"15",
16714=>X"15",
16715=>X"15",
16716=>X"15",
16717=>X"15",
16718=>X"15",
16719=>X"15",
16720=>X"15",
16721=>X"15",
16722=>X"15",
16723=>X"15",
16724=>X"15",
16725=>X"15",
16726=>X"15",
16727=>X"15",
16728=>X"15",
16729=>X"15",
16730=>X"15",
16731=>X"15",
16732=>X"15",
16733=>X"15",
16734=>X"15",
16735=>X"15",
16736=>X"15",
16737=>X"15",
16738=>X"15",
16739=>X"15",
16740=>X"00",
16741=>X"00",
16742=>X"00",
16743=>X"00",
16744=>X"00",
16745=>X"00",
16746=>X"00",
16747=>X"00",
16748=>X"00",
16749=>X"00",
16750=>X"00",
16751=>X"00",
16752=>X"00",
16753=>X"00",
16754=>X"00",
16755=>X"00",
16756=>X"00",
16757=>X"00",
16758=>X"00",
16759=>X"00",
16760=>X"00",
16761=>X"00",
16762=>X"00",
16763=>X"00",
16764=>X"00",
16765=>X"00",
16766=>X"00",
16767=>X"00",
16768=>X"00",
16769=>X"00",
16770=>X"00",
16771=>X"00",
16772=>X"00",
16773=>X"00",
16774=>X"00",
16775=>X"00",
16776=>X"00",
16777=>X"00",
16778=>X"00",
16779=>X"00",
16780=>X"00",
16781=>X"00",
16782=>X"00",
16783=>X"00",
16784=>X"00",
16785=>X"00",
16786=>X"00",
16787=>X"00",
16788=>X"00",
16789=>X"00",
16790=>X"00",
16791=>X"00",
16792=>X"00",
16793=>X"00",
16794=>X"00",
16795=>X"00",
16796=>X"00",
16797=>X"00",
16798=>X"00",
16799=>X"00",
16800=>X"00",
16801=>X"00",
16802=>X"00",
16803=>X"00",
16804=>X"00",
16805=>X"00",
16806=>X"00",
16807=>X"00",
16808=>X"00",
16809=>X"00",
16810=>X"00",
16811=>X"00",
16812=>X"00",
16813=>X"00",
16814=>X"00",
16815=>X"00",
16816=>X"00",
16817=>X"00",
16818=>X"00",
16819=>X"00",
16820=>X"00",
16821=>X"00",
16822=>X"00",
16823=>X"00",
16824=>X"00",
16825=>X"00",
16826=>X"00",
16827=>X"00",
16828=>X"00",
16829=>X"00",
16830=>X"00",
16831=>X"00",
16832=>X"00",
16833=>X"00",
16834=>X"00",
16835=>X"00",
16836=>X"00",
16837=>X"00",
16838=>X"00",
16839=>X"00",
16840=>X"00",
16841=>X"00",
16842=>X"00",
16843=>X"00",
16844=>X"00",
16845=>X"00",
16846=>X"00",
16847=>X"00",
16848=>X"00",
16849=>X"00",
16850=>X"00",
16851=>X"00",
16852=>X"00",
16853=>X"00",
16854=>X"00",
16855=>X"00",
16856=>X"00",
16857=>X"00",
16858=>X"00",
16859=>X"00",
16860=>X"00",
16861=>X"00",
16862=>X"00",
16863=>X"00",
16864=>X"00",
16865=>X"00",
16866=>X"00",
16867=>X"00",
16868=>X"00",
16869=>X"00",
16870=>X"00",
16871=>X"00",
16872=>X"00",
16873=>X"00",
16874=>X"00",
16875=>X"00",
16876=>X"00",
16877=>X"00",
16878=>X"00",
16879=>X"00",
16880=>X"00",
16881=>X"00",
16882=>X"00",
16883=>X"00",
16884=>X"00",
16885=>X"00",
16886=>X"00",
16887=>X"00",
16888=>X"00",
16889=>X"00",
16890=>X"00",
16891=>X"00",
16892=>X"00",
16893=>X"00",
16894=>X"00",
16895=>X"00",
16896=>X"04",
16897=>X"04",
16898=>X"04",
16899=>X"04",
16900=>X"04",
16901=>X"04",
16902=>X"14",
16903=>X"14",
16904=>X"14",
16905=>X"04",
16906=>X"04",
16907=>X"04",
16908=>X"15",
16909=>X"15",
16910=>X"15",
16911=>X"15",
16912=>X"15",
16913=>X"15",
16914=>X"15",
16915=>X"15",
16916=>X"15",
16917=>X"15",
16918=>X"15",
16919=>X"15",
16920=>X"29",
16921=>X"25",
16922=>X"29",
16923=>X"25",
16924=>X"25",
16925=>X"25",
16926=>X"15",
16927=>X"15",
16928=>X"15",
16929=>X"15",
16930=>X"19",
16931=>X"15",
16932=>X"19",
16933=>X"15",
16934=>X"15",
16935=>X"15",
16936=>X"15",
16937=>X"15",
16938=>X"15",
16939=>X"15",
16940=>X"15",
16941=>X"15",
16942=>X"29",
16943=>X"29",
16944=>X"3A",
16945=>X"35",
16946=>X"3A",
16947=>X"3A",
16948=>X"2A",
16949=>X"25",
16950=>X"15",
16951=>X"15",
16952=>X"15",
16953=>X"15",
16954=>X"15",
16955=>X"15",
16956=>X"15",
16957=>X"15",
16958=>X"15",
16959=>X"15",
16960=>X"15",
16961=>X"15",
16962=>X"15",
16963=>X"15",
16964=>X"15",
16965=>X"25",
16966=>X"25",
16967=>X"25",
16968=>X"25",
16969=>X"25",
16970=>X"25",
16971=>X"26",
16972=>X"36",
16973=>X"3A",
16974=>X"3B",
16975=>X"3B",
16976=>X"3F",
16977=>X"3F",
16978=>X"3F",
16979=>X"3F",
16980=>X"3F",
16981=>X"3F",
16982=>X"3F",
16983=>X"3F",
16984=>X"3F",
16985=>X"3F",
16986=>X"3F",
16987=>X"3F",
16988=>X"3F",
16989=>X"3F",
16990=>X"3F",
16991=>X"3F",
16992=>X"3F",
16993=>X"3F",
16994=>X"3F",
16995=>X"3F",
16996=>X"00",
16997=>X"00",
16998=>X"00",
16999=>X"00",
17000=>X"00",
17001=>X"00",
17002=>X"00",
17003=>X"00",
17004=>X"00",
17005=>X"00",
17006=>X"00",
17007=>X"00",
17008=>X"00",
17009=>X"00",
17010=>X"00",
17011=>X"00",
17012=>X"00",
17013=>X"00",
17014=>X"00",
17015=>X"00",
17016=>X"00",
17017=>X"00",
17018=>X"00",
17019=>X"00",
17020=>X"00",
17021=>X"00",
17022=>X"00",
17023=>X"00",
17024=>X"00",
17025=>X"00",
17026=>X"00",
17027=>X"00",
17028=>X"00",
17029=>X"00",
17030=>X"00",
17031=>X"00",
17032=>X"00",
17033=>X"00",
17034=>X"00",
17035=>X"00",
17036=>X"00",
17037=>X"00",
17038=>X"00",
17039=>X"00",
17040=>X"00",
17041=>X"00",
17042=>X"00",
17043=>X"00",
17044=>X"00",
17045=>X"00",
17046=>X"00",
17047=>X"00",
17048=>X"00",
17049=>X"00",
17050=>X"00",
17051=>X"00",
17052=>X"00",
17053=>X"00",
17054=>X"00",
17055=>X"00",
17056=>X"00",
17057=>X"00",
17058=>X"00",
17059=>X"00",
17060=>X"00",
17061=>X"00",
17062=>X"00",
17063=>X"00",
17064=>X"00",
17065=>X"00",
17066=>X"00",
17067=>X"00",
17068=>X"00",
17069=>X"00",
17070=>X"00",
17071=>X"00",
17072=>X"00",
17073=>X"00",
17074=>X"00",
17075=>X"00",
17076=>X"00",
17077=>X"00",
17078=>X"00",
17079=>X"00",
17080=>X"00",
17081=>X"00",
17082=>X"00",
17083=>X"00",
17084=>X"00",
17085=>X"00",
17086=>X"00",
17087=>X"00",
17088=>X"00",
17089=>X"00",
17090=>X"00",
17091=>X"00",
17092=>X"00",
17093=>X"00",
17094=>X"00",
17095=>X"00",
17096=>X"00",
17097=>X"00",
17098=>X"00",
17099=>X"00",
17100=>X"00",
17101=>X"00",
17102=>X"00",
17103=>X"00",
17104=>X"00",
17105=>X"00",
17106=>X"00",
17107=>X"00",
17108=>X"00",
17109=>X"00",
17110=>X"00",
17111=>X"00",
17112=>X"00",
17113=>X"00",
17114=>X"00",
17115=>X"00",
17116=>X"00",
17117=>X"00",
17118=>X"00",
17119=>X"00",
17120=>X"00",
17121=>X"00",
17122=>X"00",
17123=>X"00",
17124=>X"00",
17125=>X"00",
17126=>X"00",
17127=>X"00",
17128=>X"00",
17129=>X"00",
17130=>X"00",
17131=>X"00",
17132=>X"00",
17133=>X"00",
17134=>X"00",
17135=>X"00",
17136=>X"00",
17137=>X"00",
17138=>X"00",
17139=>X"00",
17140=>X"00",
17141=>X"00",
17142=>X"00",
17143=>X"00",
17144=>X"00",
17145=>X"00",
17146=>X"00",
17147=>X"00",
17148=>X"00",
17149=>X"00",
17150=>X"00",
17151=>X"00",
17152=>X"04",
17153=>X"04",
17154=>X"15",
17155=>X"15",
17156=>X"15",
17157=>X"15",
17158=>X"15",
17159=>X"15",
17160=>X"15",
17161=>X"15",
17162=>X"15",
17163=>X"15",
17164=>X"15",
17165=>X"15",
17166=>X"15",
17167=>X"15",
17168=>X"15",
17169=>X"15",
17170=>X"15",
17171=>X"15",
17172=>X"15",
17173=>X"15",
17174=>X"25",
17175=>X"19",
17176=>X"29",
17177=>X"2A",
17178=>X"26",
17179=>X"25",
17180=>X"2A",
17181=>X"26",
17182=>X"15",
17183=>X"15",
17184=>X"15",
17185=>X"15",
17186=>X"19",
17187=>X"15",
17188=>X"19",
17189=>X"15",
17190=>X"15",
17191=>X"15",
17192=>X"25",
17193=>X"25",
17194=>X"2A",
17195=>X"2A",
17196=>X"2A",
17197=>X"25",
17198=>X"15",
17199=>X"29",
17200=>X"2A",
17201=>X"2A",
17202=>X"3A",
17203=>X"3A",
17204=>X"3A",
17205=>X"3A",
17206=>X"2A",
17207=>X"2A",
17208=>X"2A",
17209=>X"2A",
17210=>X"3A",
17211=>X"3A",
17212=>X"3F",
17213=>X"3F",
17214=>X"3F",
17215=>X"3F",
17216=>X"3F",
17217=>X"3F",
17218=>X"3F",
17219=>X"3F",
17220=>X"3F",
17221=>X"3F",
17222=>X"3F",
17223=>X"3F",
17224=>X"3F",
17225=>X"3F",
17226=>X"3F",
17227=>X"3F",
17228=>X"3F",
17229=>X"3F",
17230=>X"3F",
17231=>X"3F",
17232=>X"3F",
17233=>X"3F",
17234=>X"3F",
17235=>X"3F",
17236=>X"3F",
17237=>X"3F",
17238=>X"3F",
17239=>X"3F",
17240=>X"3F",
17241=>X"3F",
17242=>X"3F",
17243=>X"3F",
17244=>X"3F",
17245=>X"3F",
17246=>X"3F",
17247=>X"3F",
17248=>X"3F",
17249=>X"3F",
17250=>X"3F",
17251=>X"3F",
17252=>X"00",
17253=>X"00",
17254=>X"00",
17255=>X"00",
17256=>X"00",
17257=>X"00",
17258=>X"00",
17259=>X"00",
17260=>X"00",
17261=>X"00",
17262=>X"00",
17263=>X"00",
17264=>X"00",
17265=>X"00",
17266=>X"00",
17267=>X"00",
17268=>X"00",
17269=>X"00",
17270=>X"00",
17271=>X"00",
17272=>X"00",
17273=>X"00",
17274=>X"00",
17275=>X"00",
17276=>X"00",
17277=>X"00",
17278=>X"00",
17279=>X"00",
17280=>X"00",
17281=>X"00",
17282=>X"00",
17283=>X"00",
17284=>X"00",
17285=>X"00",
17286=>X"00",
17287=>X"00",
17288=>X"00",
17289=>X"00",
17290=>X"00",
17291=>X"00",
17292=>X"00",
17293=>X"00",
17294=>X"00",
17295=>X"00",
17296=>X"00",
17297=>X"00",
17298=>X"00",
17299=>X"00",
17300=>X"00",
17301=>X"00",
17302=>X"00",
17303=>X"00",
17304=>X"00",
17305=>X"00",
17306=>X"00",
17307=>X"00",
17308=>X"00",
17309=>X"00",
17310=>X"00",
17311=>X"00",
17312=>X"00",
17313=>X"00",
17314=>X"00",
17315=>X"00",
17316=>X"00",
17317=>X"00",
17318=>X"00",
17319=>X"00",
17320=>X"00",
17321=>X"00",
17322=>X"00",
17323=>X"00",
17324=>X"00",
17325=>X"00",
17326=>X"00",
17327=>X"00",
17328=>X"00",
17329=>X"00",
17330=>X"00",
17331=>X"00",
17332=>X"00",
17333=>X"00",
17334=>X"00",
17335=>X"00",
17336=>X"00",
17337=>X"00",
17338=>X"00",
17339=>X"00",
17340=>X"00",
17341=>X"00",
17342=>X"00",
17343=>X"00",
17344=>X"00",
17345=>X"00",
17346=>X"00",
17347=>X"00",
17348=>X"00",
17349=>X"00",
17350=>X"00",
17351=>X"00",
17352=>X"00",
17353=>X"00",
17354=>X"00",
17355=>X"00",
17356=>X"00",
17357=>X"00",
17358=>X"00",
17359=>X"00",
17360=>X"00",
17361=>X"00",
17362=>X"00",
17363=>X"00",
17364=>X"00",
17365=>X"00",
17366=>X"00",
17367=>X"00",
17368=>X"00",
17369=>X"00",
17370=>X"00",
17371=>X"00",
17372=>X"00",
17373=>X"00",
17374=>X"00",
17375=>X"00",
17376=>X"00",
17377=>X"00",
17378=>X"00",
17379=>X"00",
17380=>X"00",
17381=>X"00",
17382=>X"00",
17383=>X"00",
17384=>X"00",
17385=>X"00",
17386=>X"00",
17387=>X"00",
17388=>X"00",
17389=>X"00",
17390=>X"00",
17391=>X"00",
17392=>X"00",
17393=>X"00",
17394=>X"00",
17395=>X"00",
17396=>X"00",
17397=>X"00",
17398=>X"00",
17399=>X"00",
17400=>X"00",
17401=>X"00",
17402=>X"00",
17403=>X"00",
17404=>X"00",
17405=>X"00",
17406=>X"00",
17407=>X"00",
17408=>X"15",
17409=>X"15",
17410=>X"15",
17411=>X"2A",
17412=>X"2A",
17413=>X"2A",
17414=>X"2A",
17415=>X"2A",
17416=>X"2A",
17417=>X"2A",
17418=>X"2A",
17419=>X"15",
17420=>X"15",
17421=>X"2A",
17422=>X"2A",
17423=>X"2A",
17424=>X"2A",
17425=>X"2A",
17426=>X"2E",
17427=>X"2A",
17428=>X"2A",
17429=>X"2A",
17430=>X"2B",
17431=>X"2E",
17432=>X"3A",
17433=>X"2A",
17434=>X"2B",
17435=>X"2A",
17436=>X"2A",
17437=>X"2A",
17438=>X"2A",
17439=>X"15",
17440=>X"15",
17441=>X"15",
17442=>X"15",
17443=>X"15",
17444=>X"26",
17445=>X"2A",
17446=>X"26",
17447=>X"2A",
17448=>X"2A",
17449=>X"2A",
17450=>X"2A",
17451=>X"2A",
17452=>X"2A",
17453=>X"3A",
17454=>X"2A",
17455=>X"3A",
17456=>X"3A",
17457=>X"2A",
17458=>X"3A",
17459=>X"3A",
17460=>X"3A",
17461=>X"3E",
17462=>X"3F",
17463=>X"3F",
17464=>X"3F",
17465=>X"3F",
17466=>X"3F",
17467=>X"3F",
17468=>X"3F",
17469=>X"3F",
17470=>X"3F",
17471=>X"3F",
17472=>X"3F",
17473=>X"3F",
17474=>X"3F",
17475=>X"3F",
17476=>X"3F",
17477=>X"3F",
17478=>X"3F",
17479=>X"3F",
17480=>X"3F",
17481=>X"3F",
17482=>X"3F",
17483=>X"3F",
17484=>X"3F",
17485=>X"3F",
17486=>X"3F",
17487=>X"3F",
17488=>X"3F",
17489=>X"3F",
17490=>X"3F",
17491=>X"3F",
17492=>X"3F",
17493=>X"3F",
17494=>X"3F",
17495=>X"3F",
17496=>X"3F",
17497=>X"3F",
17498=>X"3F",
17499=>X"3F",
17500=>X"3F",
17501=>X"3F",
17502=>X"3F",
17503=>X"3F",
17504=>X"3F",
17505=>X"3F",
17506=>X"3F",
17507=>X"3F",
17508=>X"00",
17509=>X"00",
17510=>X"00",
17511=>X"00",
17512=>X"00",
17513=>X"00",
17514=>X"00",
17515=>X"00",
17516=>X"00",
17517=>X"00",
17518=>X"00",
17519=>X"00",
17520=>X"00",
17521=>X"00",
17522=>X"00",
17523=>X"00",
17524=>X"00",
17525=>X"00",
17526=>X"00",
17527=>X"00",
17528=>X"00",
17529=>X"00",
17530=>X"00",
17531=>X"00",
17532=>X"00",
17533=>X"00",
17534=>X"00",
17535=>X"00",
17536=>X"00",
17537=>X"00",
17538=>X"00",
17539=>X"00",
17540=>X"00",
17541=>X"00",
17542=>X"00",
17543=>X"00",
17544=>X"00",
17545=>X"00",
17546=>X"00",
17547=>X"00",
17548=>X"00",
17549=>X"00",
17550=>X"00",
17551=>X"00",
17552=>X"00",
17553=>X"00",
17554=>X"00",
17555=>X"00",
17556=>X"00",
17557=>X"00",
17558=>X"00",
17559=>X"00",
17560=>X"00",
17561=>X"00",
17562=>X"00",
17563=>X"00",
17564=>X"00",
17565=>X"00",
17566=>X"00",
17567=>X"00",
17568=>X"00",
17569=>X"00",
17570=>X"00",
17571=>X"00",
17572=>X"00",
17573=>X"00",
17574=>X"00",
17575=>X"00",
17576=>X"00",
17577=>X"00",
17578=>X"00",
17579=>X"00",
17580=>X"00",
17581=>X"00",
17582=>X"00",
17583=>X"00",
17584=>X"00",
17585=>X"00",
17586=>X"00",
17587=>X"00",
17588=>X"00",
17589=>X"00",
17590=>X"00",
17591=>X"00",
17592=>X"00",
17593=>X"00",
17594=>X"00",
17595=>X"00",
17596=>X"00",
17597=>X"00",
17598=>X"00",
17599=>X"00",
17600=>X"00",
17601=>X"00",
17602=>X"00",
17603=>X"00",
17604=>X"00",
17605=>X"00",
17606=>X"00",
17607=>X"00",
17608=>X"00",
17609=>X"00",
17610=>X"00",
17611=>X"00",
17612=>X"00",
17613=>X"00",
17614=>X"00",
17615=>X"00",
17616=>X"00",
17617=>X"00",
17618=>X"00",
17619=>X"00",
17620=>X"00",
17621=>X"00",
17622=>X"00",
17623=>X"00",
17624=>X"00",
17625=>X"00",
17626=>X"00",
17627=>X"00",
17628=>X"00",
17629=>X"00",
17630=>X"00",
17631=>X"00",
17632=>X"00",
17633=>X"00",
17634=>X"00",
17635=>X"00",
17636=>X"00",
17637=>X"00",
17638=>X"00",
17639=>X"00",
17640=>X"00",
17641=>X"00",
17642=>X"00",
17643=>X"00",
17644=>X"00",
17645=>X"00",
17646=>X"00",
17647=>X"00",
17648=>X"00",
17649=>X"00",
17650=>X"00",
17651=>X"00",
17652=>X"00",
17653=>X"00",
17654=>X"00",
17655=>X"00",
17656=>X"00",
17657=>X"00",
17658=>X"00",
17659=>X"00",
17660=>X"00",
17661=>X"00",
17662=>X"00",
17663=>X"00",
17664=>X"3F",
17665=>X"3F",
17666=>X"3F",
17667=>X"3F",
17668=>X"3F",
17669=>X"3F",
17670=>X"3F",
17671=>X"3F",
17672=>X"3F",
17673=>X"3F",
17674=>X"3E",
17675=>X"2A",
17676=>X"2A",
17677=>X"2A",
17678=>X"3F",
17679=>X"3F",
17680=>X"3F",
17681=>X"3F",
17682=>X"3F",
17683=>X"3F",
17684=>X"3F",
17685=>X"3F",
17686=>X"3B",
17687=>X"3F",
17688=>X"3B",
17689=>X"2A",
17690=>X"2B",
17691=>X"2A",
17692=>X"2A",
17693=>X"2A",
17694=>X"2A",
17695=>X"15",
17696=>X"25",
17697=>X"25",
17698=>X"2A",
17699=>X"2A",
17700=>X"2A",
17701=>X"2A",
17702=>X"2A",
17703=>X"2A",
17704=>X"2A",
17705=>X"2A",
17706=>X"3A",
17707=>X"3A",
17708=>X"2A",
17709=>X"3A",
17710=>X"3A",
17711=>X"3A",
17712=>X"2A",
17713=>X"2A",
17714=>X"2A",
17715=>X"2A",
17716=>X"3F",
17717=>X"3F",
17718=>X"3F",
17719=>X"3F",
17720=>X"3F",
17721=>X"3F",
17722=>X"3F",
17723=>X"3F",
17724=>X"3F",
17725=>X"3F",
17726=>X"3F",
17727=>X"3F",
17728=>X"3F",
17729=>X"3F",
17730=>X"3F",
17731=>X"3F",
17732=>X"3F",
17733=>X"3F",
17734=>X"3F",
17735=>X"3F",
17736=>X"3F",
17737=>X"3F",
17738=>X"3F",
17739=>X"3F",
17740=>X"3F",
17741=>X"3F",
17742=>X"3F",
17743=>X"3F",
17744=>X"3F",
17745=>X"3F",
17746=>X"3F",
17747=>X"3F",
17748=>X"3F",
17749=>X"3F",
17750=>X"3F",
17751=>X"3F",
17752=>X"3F",
17753=>X"3F",
17754=>X"3F",
17755=>X"3E",
17756=>X"3E",
17757=>X"3F",
17758=>X"3F",
17759=>X"3F",
17760=>X"3F",
17761=>X"3F",
17762=>X"3F",
17763=>X"3F",
17764=>X"00",
17765=>X"00",
17766=>X"00",
17767=>X"00",
17768=>X"00",
17769=>X"00",
17770=>X"00",
17771=>X"00",
17772=>X"00",
17773=>X"00",
17774=>X"00",
17775=>X"00",
17776=>X"00",
17777=>X"00",
17778=>X"00",
17779=>X"00",
17780=>X"00",
17781=>X"00",
17782=>X"00",
17783=>X"00",
17784=>X"00",
17785=>X"00",
17786=>X"00",
17787=>X"00",
17788=>X"00",
17789=>X"00",
17790=>X"00",
17791=>X"00",
17792=>X"00",
17793=>X"00",
17794=>X"00",
17795=>X"00",
17796=>X"00",
17797=>X"00",
17798=>X"00",
17799=>X"00",
17800=>X"00",
17801=>X"00",
17802=>X"00",
17803=>X"00",
17804=>X"00",
17805=>X"00",
17806=>X"00",
17807=>X"00",
17808=>X"00",
17809=>X"00",
17810=>X"00",
17811=>X"00",
17812=>X"00",
17813=>X"00",
17814=>X"00",
17815=>X"00",
17816=>X"00",
17817=>X"00",
17818=>X"00",
17819=>X"00",
17820=>X"00",
17821=>X"00",
17822=>X"00",
17823=>X"00",
17824=>X"00",
17825=>X"00",
17826=>X"00",
17827=>X"00",
17828=>X"00",
17829=>X"00",
17830=>X"00",
17831=>X"00",
17832=>X"00",
17833=>X"00",
17834=>X"00",
17835=>X"00",
17836=>X"00",
17837=>X"00",
17838=>X"00",
17839=>X"00",
17840=>X"00",
17841=>X"00",
17842=>X"00",
17843=>X"00",
17844=>X"00",
17845=>X"00",
17846=>X"00",
17847=>X"00",
17848=>X"00",
17849=>X"00",
17850=>X"00",
17851=>X"00",
17852=>X"00",
17853=>X"00",
17854=>X"00",
17855=>X"00",
17856=>X"00",
17857=>X"00",
17858=>X"00",
17859=>X"00",
17860=>X"00",
17861=>X"00",
17862=>X"00",
17863=>X"00",
17864=>X"00",
17865=>X"00",
17866=>X"00",
17867=>X"00",
17868=>X"00",
17869=>X"00",
17870=>X"00",
17871=>X"00",
17872=>X"00",
17873=>X"00",
17874=>X"00",
17875=>X"00",
17876=>X"00",
17877=>X"00",
17878=>X"00",
17879=>X"00",
17880=>X"00",
17881=>X"00",
17882=>X"00",
17883=>X"00",
17884=>X"00",
17885=>X"00",
17886=>X"00",
17887=>X"00",
17888=>X"00",
17889=>X"00",
17890=>X"00",
17891=>X"00",
17892=>X"00",
17893=>X"00",
17894=>X"00",
17895=>X"00",
17896=>X"00",
17897=>X"00",
17898=>X"00",
17899=>X"00",
17900=>X"00",
17901=>X"00",
17902=>X"00",
17903=>X"00",
17904=>X"00",
17905=>X"00",
17906=>X"00",
17907=>X"00",
17908=>X"00",
17909=>X"00",
17910=>X"00",
17911=>X"00",
17912=>X"00",
17913=>X"00",
17914=>X"00",
17915=>X"00",
17916=>X"00",
17917=>X"00",
17918=>X"00",
17919=>X"00",
17920=>X"3F",
17921=>X"3F",
17922=>X"3F",
17923=>X"3F",
17924=>X"3F",
17925=>X"3F",
17926=>X"3F",
17927=>X"3F",
17928=>X"3F",
17929=>X"3F",
17930=>X"3A",
17931=>X"2A",
17932=>X"2A",
17933=>X"3F",
17934=>X"3F",
17935=>X"3F",
17936=>X"3F",
17937=>X"3A",
17938=>X"3B",
17939=>X"3B",
17940=>X"3F",
17941=>X"3F",
17942=>X"3A",
17943=>X"2A",
17944=>X"2B",
17945=>X"2A",
17946=>X"2A",
17947=>X"2A",
17948=>X"25",
17949=>X"15",
17950=>X"15",
17951=>X"25",
17952=>X"25",
17953=>X"25",
17954=>X"2A",
17955=>X"2A",
17956=>X"2A",
17957=>X"2A",
17958=>X"2A",
17959=>X"2A",
17960=>X"2A",
17961=>X"2A",
17962=>X"3A",
17963=>X"3A",
17964=>X"3A",
17965=>X"3E",
17966=>X"2A",
17967=>X"2A",
17968=>X"2A",
17969=>X"2A",
17970=>X"2A",
17971=>X"3B",
17972=>X"3F",
17973=>X"3F",
17974=>X"3F",
17975=>X"3F",
17976=>X"3F",
17977=>X"3F",
17978=>X"3F",
17979=>X"3F",
17980=>X"3F",
17981=>X"3F",
17982=>X"3F",
17983=>X"3F",
17984=>X"3F",
17985=>X"3F",
17986=>X"3F",
17987=>X"3F",
17988=>X"3F",
17989=>X"3F",
17990=>X"3F",
17991=>X"3F",
17992=>X"3F",
17993=>X"3E",
17994=>X"3F",
17995=>X"3F",
17996=>X"3F",
17997=>X"3F",
17998=>X"3F",
17999=>X"3F",
18000=>X"3F",
18001=>X"3F",
18002=>X"3F",
18003=>X"3F",
18004=>X"3F",
18005=>X"3F",
18006=>X"3F",
18007=>X"3F",
18008=>X"3F",
18009=>X"3F",
18010=>X"3F",
18011=>X"2B",
18012=>X"2A",
18013=>X"3A",
18014=>X"3E",
18015=>X"3E",
18016=>X"3A",
18017=>X"3A",
18018=>X"3A",
18019=>X"3A",
18020=>X"00",
18021=>X"00",
18022=>X"00",
18023=>X"00",
18024=>X"00",
18025=>X"00",
18026=>X"00",
18027=>X"00",
18028=>X"00",
18029=>X"00",
18030=>X"00",
18031=>X"00",
18032=>X"00",
18033=>X"00",
18034=>X"00",
18035=>X"00",
18036=>X"00",
18037=>X"00",
18038=>X"00",
18039=>X"00",
18040=>X"00",
18041=>X"00",
18042=>X"00",
18043=>X"00",
18044=>X"00",
18045=>X"00",
18046=>X"00",
18047=>X"00",
18048=>X"00",
18049=>X"00",
18050=>X"00",
18051=>X"00",
18052=>X"00",
18053=>X"00",
18054=>X"00",
18055=>X"00",
18056=>X"00",
18057=>X"00",
18058=>X"00",
18059=>X"00",
18060=>X"00",
18061=>X"00",
18062=>X"00",
18063=>X"00",
18064=>X"00",
18065=>X"00",
18066=>X"00",
18067=>X"00",
18068=>X"00",
18069=>X"00",
18070=>X"00",
18071=>X"00",
18072=>X"00",
18073=>X"00",
18074=>X"00",
18075=>X"00",
18076=>X"00",
18077=>X"00",
18078=>X"00",
18079=>X"00",
18080=>X"00",
18081=>X"00",
18082=>X"00",
18083=>X"00",
18084=>X"00",
18085=>X"00",
18086=>X"00",
18087=>X"00",
18088=>X"00",
18089=>X"00",
18090=>X"00",
18091=>X"00",
18092=>X"00",
18093=>X"00",
18094=>X"00",
18095=>X"00",
18096=>X"00",
18097=>X"00",
18098=>X"00",
18099=>X"00",
18100=>X"00",
18101=>X"00",
18102=>X"00",
18103=>X"00",
18104=>X"00",
18105=>X"00",
18106=>X"00",
18107=>X"00",
18108=>X"00",
18109=>X"00",
18110=>X"00",
18111=>X"00",
18112=>X"00",
18113=>X"00",
18114=>X"00",
18115=>X"00",
18116=>X"00",
18117=>X"00",
18118=>X"00",
18119=>X"00",
18120=>X"00",
18121=>X"00",
18122=>X"00",
18123=>X"00",
18124=>X"00",
18125=>X"00",
18126=>X"00",
18127=>X"00",
18128=>X"00",
18129=>X"00",
18130=>X"00",
18131=>X"00",
18132=>X"00",
18133=>X"00",
18134=>X"00",
18135=>X"00",
18136=>X"00",
18137=>X"00",
18138=>X"00",
18139=>X"00",
18140=>X"00",
18141=>X"00",
18142=>X"00",
18143=>X"00",
18144=>X"00",
18145=>X"00",
18146=>X"00",
18147=>X"00",
18148=>X"00",
18149=>X"00",
18150=>X"00",
18151=>X"00",
18152=>X"00",
18153=>X"00",
18154=>X"00",
18155=>X"00",
18156=>X"00",
18157=>X"00",
18158=>X"00",
18159=>X"00",
18160=>X"00",
18161=>X"00",
18162=>X"00",
18163=>X"00",
18164=>X"00",
18165=>X"00",
18166=>X"00",
18167=>X"00",
18168=>X"00",
18169=>X"00",
18170=>X"00",
18171=>X"00",
18172=>X"00",
18173=>X"00",
18174=>X"00",
18175=>X"00",
18176=>X"3F",
18177=>X"3B",
18178=>X"3F",
18179=>X"3F",
18180=>X"3F",
18181=>X"3F",
18182=>X"3F",
18183=>X"3B",
18184=>X"3A",
18185=>X"3A",
18186=>X"2A",
18187=>X"2A",
18188=>X"3F",
18189=>X"3F",
18190=>X"3F",
18191=>X"3F",
18192=>X"3F",
18193=>X"3B",
18194=>X"2F",
18195=>X"2F",
18196=>X"2A",
18197=>X"2A",
18198=>X"2A",
18199=>X"2A",
18200=>X"2A",
18201=>X"2A",
18202=>X"2A",
18203=>X"2A",
18204=>X"25",
18205=>X"2A",
18206=>X"15",
18207=>X"25",
18208=>X"29",
18209=>X"15",
18210=>X"2A",
18211=>X"2A",
18212=>X"26",
18213=>X"2A",
18214=>X"2A",
18215=>X"3A",
18216=>X"2A",
18217=>X"2A",
18218=>X"2A",
18219=>X"3F",
18220=>X"3A",
18221=>X"3A",
18222=>X"3A",
18223=>X"3E",
18224=>X"3E",
18225=>X"3A",
18226=>X"3F",
18227=>X"3B",
18228=>X"3F",
18229=>X"3F",
18230=>X"3B",
18231=>X"3B",
18232=>X"3F",
18233=>X"3F",
18234=>X"3F",
18235=>X"3F",
18236=>X"3F",
18237=>X"3F",
18238=>X"3F",
18239=>X"3E",
18240=>X"3E",
18241=>X"3F",
18242=>X"3F",
18243=>X"3E",
18244=>X"3A",
18245=>X"3A",
18246=>X"3A",
18247=>X"3F",
18248=>X"3F",
18249=>X"3F",
18250=>X"3E",
18251=>X"3F",
18252=>X"3F",
18253=>X"3F",
18254=>X"3E",
18255=>X"3A",
18256=>X"3A",
18257=>X"3B",
18258=>X"3F",
18259=>X"3F",
18260=>X"3F",
18261=>X"3F",
18262=>X"3F",
18263=>X"3F",
18264=>X"3F",
18265=>X"3F",
18266=>X"3F",
18267=>X"3F",
18268=>X"3F",
18269=>X"3F",
18270=>X"3F",
18271=>X"3F",
18272=>X"3F",
18273=>X"3A",
18274=>X"3A",
18275=>X"3A",
18276=>X"00",
18277=>X"00",
18278=>X"00",
18279=>X"00",
18280=>X"00",
18281=>X"00",
18282=>X"00",
18283=>X"00",
18284=>X"00",
18285=>X"00",
18286=>X"00",
18287=>X"00",
18288=>X"00",
18289=>X"00",
18290=>X"00",
18291=>X"00",
18292=>X"00",
18293=>X"00",
18294=>X"00",
18295=>X"00",
18296=>X"00",
18297=>X"00",
18298=>X"00",
18299=>X"00",
18300=>X"00",
18301=>X"00",
18302=>X"00",
18303=>X"00",
18304=>X"00",
18305=>X"00",
18306=>X"00",
18307=>X"00",
18308=>X"00",
18309=>X"00",
18310=>X"00",
18311=>X"00",
18312=>X"00",
18313=>X"00",
18314=>X"00",
18315=>X"00",
18316=>X"00",
18317=>X"00",
18318=>X"00",
18319=>X"00",
18320=>X"00",
18321=>X"00",
18322=>X"00",
18323=>X"00",
18324=>X"00",
18325=>X"00",
18326=>X"00",
18327=>X"00",
18328=>X"00",
18329=>X"00",
18330=>X"00",
18331=>X"00",
18332=>X"00",
18333=>X"00",
18334=>X"00",
18335=>X"00",
18336=>X"00",
18337=>X"00",
18338=>X"00",
18339=>X"00",
18340=>X"00",
18341=>X"00",
18342=>X"00",
18343=>X"00",
18344=>X"00",
18345=>X"00",
18346=>X"00",
18347=>X"00",
18348=>X"00",
18349=>X"00",
18350=>X"00",
18351=>X"00",
18352=>X"00",
18353=>X"00",
18354=>X"00",
18355=>X"00",
18356=>X"00",
18357=>X"00",
18358=>X"00",
18359=>X"00",
18360=>X"00",
18361=>X"00",
18362=>X"00",
18363=>X"00",
18364=>X"00",
18365=>X"00",
18366=>X"00",
18367=>X"00",
18368=>X"00",
18369=>X"00",
18370=>X"00",
18371=>X"00",
18372=>X"00",
18373=>X"00",
18374=>X"00",
18375=>X"00",
18376=>X"00",
18377=>X"00",
18378=>X"00",
18379=>X"00",
18380=>X"00",
18381=>X"00",
18382=>X"00",
18383=>X"00",
18384=>X"00",
18385=>X"00",
18386=>X"00",
18387=>X"00",
18388=>X"00",
18389=>X"00",
18390=>X"00",
18391=>X"00",
18392=>X"00",
18393=>X"00",
18394=>X"00",
18395=>X"00",
18396=>X"00",
18397=>X"00",
18398=>X"00",
18399=>X"00",
18400=>X"00",
18401=>X"00",
18402=>X"00",
18403=>X"00",
18404=>X"00",
18405=>X"00",
18406=>X"00",
18407=>X"00",
18408=>X"00",
18409=>X"00",
18410=>X"00",
18411=>X"00",
18412=>X"00",
18413=>X"00",
18414=>X"00",
18415=>X"00",
18416=>X"00",
18417=>X"00",
18418=>X"00",
18419=>X"00",
18420=>X"00",
18421=>X"00",
18422=>X"00",
18423=>X"00",
18424=>X"00",
18425=>X"00",
18426=>X"00",
18427=>X"00",
18428=>X"00",
18429=>X"00",
18430=>X"00",
18431=>X"00",
18432=>X"2A",
18433=>X"2A",
18434=>X"3F",
18435=>X"3A",
18436=>X"3F",
18437=>X"3B",
18438=>X"3F",
18439=>X"3F",
18440=>X"3F",
18441=>X"2A",
18442=>X"2A",
18443=>X"3F",
18444=>X"3F",
18445=>X"3F",
18446=>X"3F",
18447=>X"3B",
18448=>X"3F",
18449=>X"3B",
18450=>X"3F",
18451=>X"3F",
18452=>X"2A",
18453=>X"2A",
18454=>X"2A",
18455=>X"2A",
18456=>X"2A",
18457=>X"29",
18458=>X"15",
18459=>X"15",
18460=>X"15",
18461=>X"15",
18462=>X"15",
18463=>X"15",
18464=>X"29",
18465=>X"29",
18466=>X"2A",
18467=>X"2A",
18468=>X"2A",
18469=>X"2A",
18470=>X"2A",
18471=>X"2A",
18472=>X"2A",
18473=>X"3A",
18474=>X"3A",
18475=>X"3A",
18476=>X"3A",
18477=>X"3A",
18478=>X"3A",
18479=>X"3F",
18480=>X"3A",
18481=>X"3A",
18482=>X"3B",
18483=>X"3A",
18484=>X"3A",
18485=>X"3A",
18486=>X"3F",
18487=>X"3F",
18488=>X"3E",
18489=>X"3E",
18490=>X"3A",
18491=>X"3F",
18492=>X"3E",
18493=>X"3F",
18494=>X"3A",
18495=>X"3E",
18496=>X"3F",
18497=>X"3B",
18498=>X"3E",
18499=>X"3E",
18500=>X"3A",
18501=>X"3E",
18502=>X"3A",
18503=>X"3F",
18504=>X"3E",
18505=>X"3E",
18506=>X"3A",
18507=>X"3A",
18508=>X"3A",
18509=>X"3E",
18510=>X"3E",
18511=>X"3B",
18512=>X"3E",
18513=>X"3B",
18514=>X"3A",
18515=>X"3A",
18516=>X"3A",
18517=>X"3A",
18518=>X"3A",
18519=>X"3A",
18520=>X"3A",
18521=>X"3A",
18522=>X"3A",
18523=>X"3A",
18524=>X"3E",
18525=>X"3E",
18526=>X"3B",
18527=>X"3F",
18528=>X"3A",
18529=>X"3A",
18530=>X"3A",
18531=>X"3F",
18532=>X"00",
18533=>X"00",
18534=>X"00",
18535=>X"00",
18536=>X"00",
18537=>X"00",
18538=>X"00",
18539=>X"00",
18540=>X"00",
18541=>X"00",
18542=>X"00",
18543=>X"00",
18544=>X"00",
18545=>X"00",
18546=>X"00",
18547=>X"00",
18548=>X"00",
18549=>X"00",
18550=>X"00",
18551=>X"00",
18552=>X"00",
18553=>X"00",
18554=>X"00",
18555=>X"00",
18556=>X"00",
18557=>X"00",
18558=>X"00",
18559=>X"00",
18560=>X"00",
18561=>X"00",
18562=>X"00",
18563=>X"00",
18564=>X"00",
18565=>X"00",
18566=>X"00",
18567=>X"00",
18568=>X"00",
18569=>X"00",
18570=>X"00",
18571=>X"00",
18572=>X"00",
18573=>X"00",
18574=>X"00",
18575=>X"00",
18576=>X"00",
18577=>X"00",
18578=>X"00",
18579=>X"00",
18580=>X"00",
18581=>X"00",
18582=>X"00",
18583=>X"00",
18584=>X"00",
18585=>X"00",
18586=>X"00",
18587=>X"00",
18588=>X"00",
18589=>X"00",
18590=>X"00",
18591=>X"00",
18592=>X"00",
18593=>X"00",
18594=>X"00",
18595=>X"00",
18596=>X"00",
18597=>X"00",
18598=>X"00",
18599=>X"00",
18600=>X"00",
18601=>X"00",
18602=>X"00",
18603=>X"00",
18604=>X"00",
18605=>X"00",
18606=>X"00",
18607=>X"00",
18608=>X"00",
18609=>X"00",
18610=>X"00",
18611=>X"00",
18612=>X"00",
18613=>X"00",
18614=>X"00",
18615=>X"00",
18616=>X"00",
18617=>X"00",
18618=>X"00",
18619=>X"00",
18620=>X"00",
18621=>X"00",
18622=>X"00",
18623=>X"00",
18624=>X"00",
18625=>X"00",
18626=>X"00",
18627=>X"00",
18628=>X"00",
18629=>X"00",
18630=>X"00",
18631=>X"00",
18632=>X"00",
18633=>X"00",
18634=>X"00",
18635=>X"00",
18636=>X"00",
18637=>X"00",
18638=>X"00",
18639=>X"00",
18640=>X"00",
18641=>X"00",
18642=>X"00",
18643=>X"00",
18644=>X"00",
18645=>X"00",
18646=>X"00",
18647=>X"00",
18648=>X"00",
18649=>X"00",
18650=>X"00",
18651=>X"00",
18652=>X"00",
18653=>X"00",
18654=>X"00",
18655=>X"00",
18656=>X"00",
18657=>X"00",
18658=>X"00",
18659=>X"00",
18660=>X"00",
18661=>X"00",
18662=>X"00",
18663=>X"00",
18664=>X"00",
18665=>X"00",
18666=>X"00",
18667=>X"00",
18668=>X"00",
18669=>X"00",
18670=>X"00",
18671=>X"00",
18672=>X"00",
18673=>X"00",
18674=>X"00",
18675=>X"00",
18676=>X"00",
18677=>X"00",
18678=>X"00",
18679=>X"00",
18680=>X"00",
18681=>X"00",
18682=>X"00",
18683=>X"00",
18684=>X"00",
18685=>X"00",
18686=>X"00",
18687=>X"00",
18688=>X"2A",
18689=>X"2A",
18690=>X"2A",
18691=>X"3A",
18692=>X"3A",
18693=>X"3A",
18694=>X"3A",
18695=>X"2A",
18696=>X"2A",
18697=>X"26",
18698=>X"2A",
18699=>X"3F",
18700=>X"3E",
18701=>X"2A",
18702=>X"2A",
18703=>X"3A",
18704=>X"3A",
18705=>X"2A",
18706=>X"2A",
18707=>X"2A",
18708=>X"2A",
18709=>X"2A",
18710=>X"2A",
18711=>X"26",
18712=>X"26",
18713=>X"26",
18714=>X"15",
18715=>X"25",
18716=>X"26",
18717=>X"25",
18718=>X"25",
18719=>X"15",
18720=>X"25",
18721=>X"26",
18722=>X"25",
18723=>X"2A",
18724=>X"29",
18725=>X"2A",
18726=>X"2A",
18727=>X"29",
18728=>X"29",
18729=>X"3A",
18730=>X"3A",
18731=>X"2A",
18732=>X"2A",
18733=>X"3A",
18734=>X"3A",
18735=>X"2A",
18736=>X"3A",
18737=>X"2A",
18738=>X"2A",
18739=>X"3A",
18740=>X"3A",
18741=>X"3A",
18742=>X"3E",
18743=>X"3A",
18744=>X"3A",
18745=>X"3E",
18746=>X"3A",
18747=>X"3A",
18748=>X"3A",
18749=>X"3A",
18750=>X"3A",
18751=>X"3A",
18752=>X"3A",
18753=>X"3A",
18754=>X"3A",
18755=>X"3E",
18756=>X"3A",
18757=>X"3A",
18758=>X"3A",
18759=>X"3A",
18760=>X"3A",
18761=>X"3A",
18762=>X"3A",
18763=>X"3A",
18764=>X"3A",
18765=>X"3E",
18766=>X"3E",
18767=>X"2A",
18768=>X"3A",
18769=>X"3A",
18770=>X"3A",
18771=>X"3A",
18772=>X"2A",
18773=>X"2A",
18774=>X"2A",
18775=>X"2A",
18776=>X"2A",
18777=>X"2A",
18778=>X"2A",
18779=>X"2A",
18780=>X"2A",
18781=>X"2A",
18782=>X"2A",
18783=>X"2A",
18784=>X"2A",
18785=>X"2A",
18786=>X"3A",
18787=>X"2A",
18788=>X"00",
18789=>X"00",
18790=>X"00",
18791=>X"00",
18792=>X"00",
18793=>X"00",
18794=>X"00",
18795=>X"00",
18796=>X"00",
18797=>X"00",
18798=>X"00",
18799=>X"00",
18800=>X"00",
18801=>X"00",
18802=>X"00",
18803=>X"00",
18804=>X"00",
18805=>X"00",
18806=>X"00",
18807=>X"00",
18808=>X"00",
18809=>X"00",
18810=>X"00",
18811=>X"00",
18812=>X"00",
18813=>X"00",
18814=>X"00",
18815=>X"00",
18816=>X"00",
18817=>X"00",
18818=>X"00",
18819=>X"00",
18820=>X"00",
18821=>X"00",
18822=>X"00",
18823=>X"00",
18824=>X"00",
18825=>X"00",
18826=>X"00",
18827=>X"00",
18828=>X"00",
18829=>X"00",
18830=>X"00",
18831=>X"00",
18832=>X"00",
18833=>X"00",
18834=>X"00",
18835=>X"00",
18836=>X"00",
18837=>X"00",
18838=>X"00",
18839=>X"00",
18840=>X"00",
18841=>X"00",
18842=>X"00",
18843=>X"00",
18844=>X"00",
18845=>X"00",
18846=>X"00",
18847=>X"00",
18848=>X"00",
18849=>X"00",
18850=>X"00",
18851=>X"00",
18852=>X"00",
18853=>X"00",
18854=>X"00",
18855=>X"00",
18856=>X"00",
18857=>X"00",
18858=>X"00",
18859=>X"00",
18860=>X"00",
18861=>X"00",
18862=>X"00",
18863=>X"00",
18864=>X"00",
18865=>X"00",
18866=>X"00",
18867=>X"00",
18868=>X"00",
18869=>X"00",
18870=>X"00",
18871=>X"00",
18872=>X"00",
18873=>X"00",
18874=>X"00",
18875=>X"00",
18876=>X"00",
18877=>X"00",
18878=>X"00",
18879=>X"00",
18880=>X"00",
18881=>X"00",
18882=>X"00",
18883=>X"00",
18884=>X"00",
18885=>X"00",
18886=>X"00",
18887=>X"00",
18888=>X"00",
18889=>X"00",
18890=>X"00",
18891=>X"00",
18892=>X"00",
18893=>X"00",
18894=>X"00",
18895=>X"00",
18896=>X"00",
18897=>X"00",
18898=>X"00",
18899=>X"00",
18900=>X"00",
18901=>X"00",
18902=>X"00",
18903=>X"00",
18904=>X"00",
18905=>X"00",
18906=>X"00",
18907=>X"00",
18908=>X"00",
18909=>X"00",
18910=>X"00",
18911=>X"00",
18912=>X"00",
18913=>X"00",
18914=>X"00",
18915=>X"00",
18916=>X"00",
18917=>X"00",
18918=>X"00",
18919=>X"00",
18920=>X"00",
18921=>X"00",
18922=>X"00",
18923=>X"00",
18924=>X"00",
18925=>X"00",
18926=>X"00",
18927=>X"00",
18928=>X"00",
18929=>X"00",
18930=>X"00",
18931=>X"00",
18932=>X"00",
18933=>X"00",
18934=>X"00",
18935=>X"00",
18936=>X"00",
18937=>X"00",
18938=>X"00",
18939=>X"00",
18940=>X"00",
18941=>X"00",
18942=>X"00",
18943=>X"00",
18944=>X"2A",
18945=>X"2A",
18946=>X"2A",
18947=>X"2A",
18948=>X"2A",
18949=>X"2A",
18950=>X"2A",
18951=>X"2A",
18952=>X"26",
18953=>X"26",
18954=>X"2A",
18955=>X"2A",
18956=>X"2A",
18957=>X"2A",
18958=>X"2A",
18959=>X"2A",
18960=>X"2A",
18961=>X"2A",
18962=>X"25",
18963=>X"25",
18964=>X"25",
18965=>X"25",
18966=>X"15",
18967=>X"15",
18968=>X"2A",
18969=>X"26",
18970=>X"15",
18971=>X"15",
18972=>X"25",
18973=>X"25",
18974=>X"15",
18975=>X"15",
18976=>X"25",
18977=>X"29",
18978=>X"25",
18979=>X"25",
18980=>X"29",
18981=>X"29",
18982=>X"25",
18983=>X"25",
18984=>X"25",
18985=>X"25",
18986=>X"2A",
18987=>X"2A",
18988=>X"2A",
18989=>X"2A",
18990=>X"2A",
18991=>X"2A",
18992=>X"2A",
18993=>X"2A",
18994=>X"2A",
18995=>X"2A",
18996=>X"2A",
18997=>X"2A",
18998=>X"2A",
18999=>X"2A",
19000=>X"2A",
19001=>X"2A",
19002=>X"2A",
19003=>X"2A",
19004=>X"2A",
19005=>X"2A",
19006=>X"2A",
19007=>X"2A",
19008=>X"2A",
19009=>X"2A",
19010=>X"3A",
19011=>X"3A",
19012=>X"3A",
19013=>X"3A",
19014=>X"3A",
19015=>X"3A",
19016=>X"2A",
19017=>X"2A",
19018=>X"3A",
19019=>X"3A",
19020=>X"2A",
19021=>X"2A",
19022=>X"2A",
19023=>X"2A",
19024=>X"29",
19025=>X"29",
19026=>X"29",
19027=>X"29",
19028=>X"29",
19029=>X"29",
19030=>X"25",
19031=>X"25",
19032=>X"25",
19033=>X"25",
19034=>X"25",
19035=>X"25",
19036=>X"25",
19037=>X"25",
19038=>X"29",
19039=>X"29",
19040=>X"2A",
19041=>X"2A",
19042=>X"25",
19043=>X"25",
19044=>X"00",
19045=>X"00",
19046=>X"00",
19047=>X"00",
19048=>X"00",
19049=>X"00",
19050=>X"00",
19051=>X"00",
19052=>X"00",
19053=>X"00",
19054=>X"00",
19055=>X"00",
19056=>X"00",
19057=>X"00",
19058=>X"00",
19059=>X"00",
19060=>X"00",
19061=>X"00",
19062=>X"00",
19063=>X"00",
19064=>X"00",
19065=>X"00",
19066=>X"00",
19067=>X"00",
19068=>X"00",
19069=>X"00",
19070=>X"00",
19071=>X"00",
19072=>X"00",
19073=>X"00",
19074=>X"00",
19075=>X"00",
19076=>X"00",
19077=>X"00",
19078=>X"00",
19079=>X"00",
19080=>X"00",
19081=>X"00",
19082=>X"00",
19083=>X"00",
19084=>X"00",
19085=>X"00",
19086=>X"00",
19087=>X"00",
19088=>X"00",
19089=>X"00",
19090=>X"00",
19091=>X"00",
19092=>X"00",
19093=>X"00",
19094=>X"00",
19095=>X"00",
19096=>X"00",
19097=>X"00",
19098=>X"00",
19099=>X"00",
19100=>X"00",
19101=>X"00",
19102=>X"00",
19103=>X"00",
19104=>X"00",
19105=>X"00",
19106=>X"00",
19107=>X"00",
19108=>X"00",
19109=>X"00",
19110=>X"00",
19111=>X"00",
19112=>X"00",
19113=>X"00",
19114=>X"00",
19115=>X"00",
19116=>X"00",
19117=>X"00",
19118=>X"00",
19119=>X"00",
19120=>X"00",
19121=>X"00",
19122=>X"00",
19123=>X"00",
19124=>X"00",
19125=>X"00",
19126=>X"00",
19127=>X"00",
19128=>X"00",
19129=>X"00",
19130=>X"00",
19131=>X"00",
19132=>X"00",
19133=>X"00",
19134=>X"00",
19135=>X"00",
19136=>X"00",
19137=>X"00",
19138=>X"00",
19139=>X"00",
19140=>X"00",
19141=>X"00",
19142=>X"00",
19143=>X"00",
19144=>X"00",
19145=>X"00",
19146=>X"00",
19147=>X"00",
19148=>X"00",
19149=>X"00",
19150=>X"00",
19151=>X"00",
19152=>X"00",
19153=>X"00",
19154=>X"00",
19155=>X"00",
19156=>X"00",
19157=>X"00",
19158=>X"00",
19159=>X"00",
19160=>X"00",
19161=>X"00",
19162=>X"00",
19163=>X"00",
19164=>X"00",
19165=>X"00",
19166=>X"00",
19167=>X"00",
19168=>X"00",
19169=>X"00",
19170=>X"00",
19171=>X"00",
19172=>X"00",
19173=>X"00",
19174=>X"00",
19175=>X"00",
19176=>X"00",
19177=>X"00",
19178=>X"00",
19179=>X"00",
19180=>X"00",
19181=>X"00",
19182=>X"00",
19183=>X"00",
19184=>X"00",
19185=>X"00",
19186=>X"00",
19187=>X"00",
19188=>X"00",
19189=>X"00",
19190=>X"00",
19191=>X"00",
19192=>X"00",
19193=>X"00",
19194=>X"00",
19195=>X"00",
19196=>X"00",
19197=>X"00",
19198=>X"00",
19199=>X"00",
19200=>X"00",
19201=>X"00",
19202=>X"00",
19203=>X"00",
19204=>X"00",
19205=>X"00",
19206=>X"00",
19207=>X"00",
19208=>X"00",
19209=>X"00",
19210=>X"00",
19211=>X"00",
19212=>X"00",
19213=>X"00",
19214=>X"00",
19215=>X"00",
19216=>X"00",
19217=>X"00",
19218=>X"00",
19219=>X"00",
19220=>X"00",
19221=>X"00",
19222=>X"00",
19223=>X"00",
19224=>X"00",
19225=>X"00",
19226=>X"00",
19227=>X"00",
19228=>X"00",
19229=>X"00",
19230=>X"00",
19231=>X"00",
19232=>X"00",
19233=>X"00",
19234=>X"00",
19235=>X"00",
19236=>X"00",
19237=>X"00",
19238=>X"00",
19239=>X"00",
19240=>X"00",
19241=>X"00",
19242=>X"00",
19243=>X"00",
19244=>X"00",
19245=>X"00",
19246=>X"00",
19247=>X"00",
19248=>X"00",
19249=>X"00",
19250=>X"00",
19251=>X"00",
19252=>X"00",
19253=>X"00",
19254=>X"00",
19255=>X"00",
19256=>X"00",
19257=>X"00",
19258=>X"00",
19259=>X"00",
19260=>X"00",
19261=>X"00",
19262=>X"00",
19263=>X"00",
19264=>X"00",
19265=>X"00",
19266=>X"00",
19267=>X"00",
19268=>X"00",
19269=>X"00",
19270=>X"00",
19271=>X"00",
19272=>X"00",
19273=>X"00",
19274=>X"00",
19275=>X"00",
19276=>X"00",
19277=>X"00",
19278=>X"00",
19279=>X"00",
19280=>X"00",
19281=>X"00",
19282=>X"00",
19283=>X"00",
19284=>X"00",
19285=>X"00",
19286=>X"00",
19287=>X"00",
19288=>X"00",
19289=>X"00",
19290=>X"00",
19291=>X"00",
19292=>X"00",
19293=>X"00",
19294=>X"00",
19295=>X"00",
19296=>X"00",
19297=>X"00",
19298=>X"00",
19299=>X"00",
19300=>X"00",
19301=>X"00",
19302=>X"00",
19303=>X"00",
19304=>X"00",
19305=>X"00",
19306=>X"00",
19307=>X"00",
19308=>X"00",
19309=>X"00",
19310=>X"00",
19311=>X"00",
19312=>X"00",
19313=>X"00",
19314=>X"00",
19315=>X"00",
19316=>X"00",
19317=>X"00",
19318=>X"00",
19319=>X"00",
19320=>X"00",
19321=>X"00",
19322=>X"00",
19323=>X"00",
19324=>X"00",
19325=>X"00",
19326=>X"00",
19327=>X"00",
19328=>X"00",
19329=>X"00",
19330=>X"00",
19331=>X"00",
19332=>X"00",
19333=>X"00",
19334=>X"00",
19335=>X"00",
19336=>X"00",
19337=>X"00",
19338=>X"00",
19339=>X"00",
19340=>X"00",
19341=>X"00",
19342=>X"00",
19343=>X"00",
19344=>X"00",
19345=>X"00",
19346=>X"00",
19347=>X"00",
19348=>X"00",
19349=>X"00",
19350=>X"00",
19351=>X"00",
19352=>X"00",
19353=>X"00",
19354=>X"00",
19355=>X"00",
19356=>X"00",
19357=>X"00",
19358=>X"00",
19359=>X"00",
19360=>X"00",
19361=>X"00",
19362=>X"00",
19363=>X"00",
19364=>X"00",
19365=>X"00",
19366=>X"00",
19367=>X"00",
19368=>X"00",
19369=>X"00",
19370=>X"00",
19371=>X"00",
19372=>X"00",
19373=>X"00",
19374=>X"00",
19375=>X"00",
19376=>X"00",
19377=>X"00",
19378=>X"00",
19379=>X"00",
19380=>X"00",
19381=>X"00",
19382=>X"00",
19383=>X"00",
19384=>X"00",
19385=>X"00",
19386=>X"00",
19387=>X"00",
19388=>X"00",
19389=>X"00",
19390=>X"00",
19391=>X"00",
19392=>X"00",
19393=>X"00",
19394=>X"00",
19395=>X"00",
19396=>X"00",
19397=>X"00",
19398=>X"00",
19399=>X"00",
19400=>X"00",
19401=>X"00",
19402=>X"00",
19403=>X"00",
19404=>X"00",
19405=>X"00",
19406=>X"00",
19407=>X"00",
19408=>X"00",
19409=>X"00",
19410=>X"00",
19411=>X"00",
19412=>X"00",
19413=>X"00",
19414=>X"00",
19415=>X"00",
19416=>X"00",
19417=>X"00",
19418=>X"00",
19419=>X"00",
19420=>X"00",
19421=>X"00",
19422=>X"00",
19423=>X"00",
19424=>X"00",
19425=>X"00",
19426=>X"00",
19427=>X"00",
19428=>X"00",
19429=>X"00",
19430=>X"00",
19431=>X"00",
19432=>X"00",
19433=>X"00",
19434=>X"00",
19435=>X"00",
19436=>X"00",
19437=>X"00",
19438=>X"00",
19439=>X"00",
19440=>X"00",
19441=>X"00",
19442=>X"00",
19443=>X"00",
19444=>X"00",
19445=>X"00",
19446=>X"00",
19447=>X"00",
19448=>X"00",
19449=>X"00",
19450=>X"00",
19451=>X"00",
19452=>X"00",
19453=>X"00",
19454=>X"00",
19455=>X"00",
19456=>X"00",
19457=>X"00",
19458=>X"00",
19459=>X"00",
19460=>X"00",
19461=>X"00",
19462=>X"00",
19463=>X"00",
19464=>X"00",
19465=>X"00",
19466=>X"00",
19467=>X"00",
19468=>X"00",
19469=>X"00",
19470=>X"00",
19471=>X"00",
19472=>X"00",
19473=>X"00",
19474=>X"00",
19475=>X"00",
19476=>X"00",
19477=>X"00",
19478=>X"00",
19479=>X"00",
19480=>X"00",
19481=>X"00",
19482=>X"00",
19483=>X"00",
19484=>X"00",
19485=>X"00",
19486=>X"00",
19487=>X"00",
19488=>X"00",
19489=>X"00",
19490=>X"00",
19491=>X"00",
19492=>X"00",
19493=>X"00",
19494=>X"00",
19495=>X"00",
19496=>X"00",
19497=>X"00",
19498=>X"00",
19499=>X"00",
19500=>X"00",
19501=>X"00",
19502=>X"00",
19503=>X"00",
19504=>X"00",
19505=>X"00",
19506=>X"00",
19507=>X"00",
19508=>X"00",
19509=>X"00",
19510=>X"00",
19511=>X"00",
19512=>X"00",
19513=>X"00",
19514=>X"00",
19515=>X"00",
19516=>X"00",
19517=>X"00",
19518=>X"00",
19519=>X"00",
19520=>X"00",
19521=>X"00",
19522=>X"00",
19523=>X"00",
19524=>X"00",
19525=>X"00",
19526=>X"00",
19527=>X"00",
19528=>X"00",
19529=>X"00",
19530=>X"00",
19531=>X"00",
19532=>X"00",
19533=>X"00",
19534=>X"00",
19535=>X"00",
19536=>X"00",
19537=>X"00",
19538=>X"00",
19539=>X"00",
19540=>X"00",
19541=>X"00",
19542=>X"00",
19543=>X"00",
19544=>X"00",
19545=>X"00",
19546=>X"00",
19547=>X"00",
19548=>X"00",
19549=>X"00",
19550=>X"00",
19551=>X"00",
19552=>X"00",
19553=>X"00",
19554=>X"00",
19555=>X"00",
19556=>X"00",
19557=>X"00",
19558=>X"00",
19559=>X"00",
19560=>X"00",
19561=>X"00",
19562=>X"00",
19563=>X"00",
19564=>X"00",
19565=>X"00",
19566=>X"00",
19567=>X"00",
19568=>X"00",
19569=>X"00",
19570=>X"00",
19571=>X"00",
19572=>X"00",
19573=>X"00",
19574=>X"00",
19575=>X"00",
19576=>X"00",
19577=>X"00",
19578=>X"00",
19579=>X"00",
19580=>X"00",
19581=>X"00",
19582=>X"00",
19583=>X"00",
19584=>X"00",
19585=>X"00",
19586=>X"00",
19587=>X"00",
19588=>X"00",
19589=>X"00",
19590=>X"00",
19591=>X"00",
19592=>X"00",
19593=>X"00",
19594=>X"00",
19595=>X"00",
19596=>X"00",
19597=>X"00",
19598=>X"00",
19599=>X"00",
19600=>X"00",
19601=>X"00",
19602=>X"00",
19603=>X"00",
19604=>X"00",
19605=>X"00",
19606=>X"00",
19607=>X"00",
19608=>X"00",
19609=>X"00",
19610=>X"00",
19611=>X"00",
19612=>X"00",
19613=>X"00",
19614=>X"00",
19615=>X"00",
19616=>X"00",
19617=>X"00",
19618=>X"00",
19619=>X"00",
19620=>X"00",
19621=>X"00",
19622=>X"00",
19623=>X"00",
19624=>X"00",
19625=>X"00",
19626=>X"00",
19627=>X"00",
19628=>X"00",
19629=>X"00",
19630=>X"00",
19631=>X"00",
19632=>X"00",
19633=>X"00",
19634=>X"00",
19635=>X"00",
19636=>X"00",
19637=>X"00",
19638=>X"00",
19639=>X"00",
19640=>X"00",
19641=>X"00",
19642=>X"00",
19643=>X"00",
19644=>X"00",
19645=>X"00",
19646=>X"00",
19647=>X"00",
19648=>X"00",
19649=>X"00",
19650=>X"00",
19651=>X"00",
19652=>X"00",
19653=>X"00",
19654=>X"00",
19655=>X"00",
19656=>X"00",
19657=>X"00",
19658=>X"00",
19659=>X"00",
19660=>X"00",
19661=>X"00",
19662=>X"00",
19663=>X"00",
19664=>X"00",
19665=>X"00",
19666=>X"00",
19667=>X"00",
19668=>X"00",
19669=>X"00",
19670=>X"00",
19671=>X"00",
19672=>X"00",
19673=>X"00",
19674=>X"00",
19675=>X"00",
19676=>X"00",
19677=>X"00",
19678=>X"00",
19679=>X"00",
19680=>X"00",
19681=>X"00",
19682=>X"00",
19683=>X"00",
19684=>X"00",
19685=>X"00",
19686=>X"00",
19687=>X"00",
19688=>X"00",
19689=>X"00",
19690=>X"00",
19691=>X"00",
19692=>X"00",
19693=>X"00",
19694=>X"00",
19695=>X"00",
19696=>X"00",
19697=>X"00",
19698=>X"00",
19699=>X"00",
19700=>X"00",
19701=>X"00",
19702=>X"00",
19703=>X"00",
19704=>X"00",
19705=>X"00",
19706=>X"00",
19707=>X"00",
19708=>X"00",
19709=>X"00",
19710=>X"00",
19711=>X"00",
19712=>X"00",
19713=>X"00",
19714=>X"00",
19715=>X"00",
19716=>X"00",
19717=>X"00",
19718=>X"00",
19719=>X"00",
19720=>X"00",
19721=>X"00",
19722=>X"00",
19723=>X"00",
19724=>X"00",
19725=>X"00",
19726=>X"00",
19727=>X"00",
19728=>X"00",
19729=>X"00",
19730=>X"00",
19731=>X"00",
19732=>X"00",
19733=>X"00",
19734=>X"00",
19735=>X"00",
19736=>X"00",
19737=>X"00",
19738=>X"00",
19739=>X"00",
19740=>X"00",
19741=>X"00",
19742=>X"00",
19743=>X"00",
19744=>X"00",
19745=>X"00",
19746=>X"00",
19747=>X"00",
19748=>X"00",
19749=>X"00",
19750=>X"00",
19751=>X"00",
19752=>X"00",
19753=>X"00",
19754=>X"00",
19755=>X"00",
19756=>X"00",
19757=>X"00",
19758=>X"00",
19759=>X"00",
19760=>X"00",
19761=>X"00",
19762=>X"00",
19763=>X"00",
19764=>X"00",
19765=>X"00",
19766=>X"00",
19767=>X"00",
19768=>X"00",
19769=>X"00",
19770=>X"00",
19771=>X"00",
19772=>X"00",
19773=>X"00",
19774=>X"00",
19775=>X"00",
19776=>X"00",
19777=>X"00",
19778=>X"00",
19779=>X"00",
19780=>X"00",
19781=>X"00",
19782=>X"00",
19783=>X"00",
19784=>X"00",
19785=>X"00",
19786=>X"00",
19787=>X"00",
19788=>X"00",
19789=>X"00",
19790=>X"00",
19791=>X"00",
19792=>X"00",
19793=>X"00",
19794=>X"00",
19795=>X"00",
19796=>X"00",
19797=>X"00",
19798=>X"00",
19799=>X"00",
19800=>X"00",
19801=>X"00",
19802=>X"00",
19803=>X"00",
19804=>X"00",
19805=>X"00",
19806=>X"00",
19807=>X"00",
19808=>X"00",
19809=>X"00",
19810=>X"00",
19811=>X"00",
19812=>X"00",
19813=>X"00",
19814=>X"00",
19815=>X"00",
19816=>X"00",
19817=>X"00",
19818=>X"00",
19819=>X"00",
19820=>X"00",
19821=>X"00",
19822=>X"00",
19823=>X"00",
19824=>X"00",
19825=>X"00",
19826=>X"00",
19827=>X"00",
19828=>X"00",
19829=>X"00",
19830=>X"00",
19831=>X"00",
19832=>X"00",
19833=>X"00",
19834=>X"00",
19835=>X"00",
19836=>X"00",
19837=>X"00",
19838=>X"00",
19839=>X"00",
19840=>X"00",
19841=>X"00",
19842=>X"00",
19843=>X"00",
19844=>X"00",
19845=>X"00",
19846=>X"00",
19847=>X"00",
19848=>X"00",
19849=>X"00",
19850=>X"00",
19851=>X"00",
19852=>X"00",
19853=>X"00",
19854=>X"00",
19855=>X"00",
19856=>X"00",
19857=>X"00",
19858=>X"00",
19859=>X"00",
19860=>X"00",
19861=>X"00",
19862=>X"00",
19863=>X"00",
19864=>X"00",
19865=>X"00",
19866=>X"00",
19867=>X"00",
19868=>X"00",
19869=>X"00",
19870=>X"00",
19871=>X"00",
19872=>X"00",
19873=>X"00",
19874=>X"00",
19875=>X"00",
19876=>X"00",
19877=>X"00",
19878=>X"00",
19879=>X"00",
19880=>X"00",
19881=>X"00",
19882=>X"00",
19883=>X"00",
19884=>X"00",
19885=>X"00",
19886=>X"00",
19887=>X"00",
19888=>X"00",
19889=>X"00",
19890=>X"00",
19891=>X"00",
19892=>X"00",
19893=>X"00",
19894=>X"00",
19895=>X"00",
19896=>X"00",
19897=>X"00",
19898=>X"00",
19899=>X"00",
19900=>X"00",
19901=>X"00",
19902=>X"00",
19903=>X"00",
19904=>X"00",
19905=>X"00",
19906=>X"00",
19907=>X"00",
19908=>X"00",
19909=>X"00",
19910=>X"00",
19911=>X"00",
19912=>X"00",
19913=>X"00",
19914=>X"00",
19915=>X"00",
19916=>X"00",
19917=>X"00",
19918=>X"00",
19919=>X"00",
19920=>X"00",
19921=>X"00",
19922=>X"00",
19923=>X"00",
19924=>X"00",
19925=>X"00",
19926=>X"00",
19927=>X"00",
19928=>X"00",
19929=>X"00",
19930=>X"00",
19931=>X"00",
19932=>X"00",
19933=>X"00",
19934=>X"00",
19935=>X"00",
19936=>X"00",
19937=>X"00",
19938=>X"00",
19939=>X"00",
19940=>X"00",
19941=>X"00",
19942=>X"00",
19943=>X"00",
19944=>X"00",
19945=>X"00",
19946=>X"00",
19947=>X"00",
19948=>X"00",
19949=>X"00",
19950=>X"00",
19951=>X"00",
19952=>X"00",
19953=>X"00",
19954=>X"00",
19955=>X"00",
19956=>X"00",
19957=>X"00",
19958=>X"00",
19959=>X"00",
19960=>X"00",
19961=>X"00",
19962=>X"00",
19963=>X"00",
19964=>X"00",
19965=>X"00",
19966=>X"00",
19967=>X"00",
19968=>X"00",
19969=>X"00",
19970=>X"00",
19971=>X"00",
19972=>X"00",
19973=>X"00",
19974=>X"00",
19975=>X"00",
19976=>X"00",
19977=>X"00",
19978=>X"00",
19979=>X"00",
19980=>X"00",
19981=>X"00",
19982=>X"00",
19983=>X"00",
19984=>X"00",
19985=>X"00",
19986=>X"00",
19987=>X"00",
19988=>X"00",
19989=>X"00",
19990=>X"00",
19991=>X"00",
19992=>X"00",
19993=>X"00",
19994=>X"00",
19995=>X"00",
19996=>X"00",
19997=>X"00",
19998=>X"00",
19999=>X"00",
20000=>X"00",
20001=>X"00",
20002=>X"00",
20003=>X"00",
20004=>X"00",
20005=>X"00",
20006=>X"00",
20007=>X"00",
20008=>X"00",
20009=>X"00",
20010=>X"00",
20011=>X"00",
20012=>X"00",
20013=>X"00",
20014=>X"00",
20015=>X"00",
20016=>X"00",
20017=>X"00",
20018=>X"00",
20019=>X"00",
20020=>X"00",
20021=>X"00",
20022=>X"00",
20023=>X"00",
20024=>X"00",
20025=>X"00",
20026=>X"00",
20027=>X"00",
20028=>X"00",
20029=>X"00",
20030=>X"00",
20031=>X"00",
20032=>X"00",
20033=>X"00",
20034=>X"00",
20035=>X"00",
20036=>X"00",
20037=>X"00",
20038=>X"00",
20039=>X"00",
20040=>X"00",
20041=>X"00",
20042=>X"00",
20043=>X"00",
20044=>X"00",
20045=>X"00",
20046=>X"00",
20047=>X"00",
20048=>X"00",
20049=>X"00",
20050=>X"00",
20051=>X"00",
20052=>X"00",
20053=>X"00",
20054=>X"00",
20055=>X"00",
20056=>X"00",
20057=>X"00",
20058=>X"00",
20059=>X"00",
20060=>X"00",
20061=>X"00",
20062=>X"00",
20063=>X"00",
20064=>X"00",
20065=>X"00",
20066=>X"00",
20067=>X"00",
20068=>X"00",
20069=>X"00",
20070=>X"00",
20071=>X"00",
20072=>X"00",
20073=>X"00",
20074=>X"00",
20075=>X"00",
20076=>X"00",
20077=>X"00",
20078=>X"00",
20079=>X"00",
20080=>X"00",
20081=>X"00",
20082=>X"00",
20083=>X"00",
20084=>X"00",
20085=>X"00",
20086=>X"00",
20087=>X"00",
20088=>X"00",
20089=>X"00",
20090=>X"00",
20091=>X"00",
20092=>X"00",
20093=>X"00",
20094=>X"00",
20095=>X"00",
20096=>X"00",
20097=>X"00",
20098=>X"00",
20099=>X"00",
20100=>X"00",
20101=>X"00",
20102=>X"00",
20103=>X"00",
20104=>X"00",
20105=>X"00",
20106=>X"00",
20107=>X"00",
20108=>X"00",
20109=>X"00",
20110=>X"00",
20111=>X"00",
20112=>X"00",
20113=>X"00",
20114=>X"00",
20115=>X"00",
20116=>X"00",
20117=>X"00",
20118=>X"00",
20119=>X"00",
20120=>X"00",
20121=>X"00",
20122=>X"00",
20123=>X"00",
20124=>X"00",
20125=>X"00",
20126=>X"00",
20127=>X"00",
20128=>X"00",
20129=>X"00",
20130=>X"00",
20131=>X"00",
20132=>X"00",
20133=>X"00",
20134=>X"00",
20135=>X"00",
20136=>X"00",
20137=>X"00",
20138=>X"00",
20139=>X"00",
20140=>X"00",
20141=>X"00",
20142=>X"00",
20143=>X"00",
20144=>X"00",
20145=>X"00",
20146=>X"00",
20147=>X"00",
20148=>X"00",
20149=>X"00",
20150=>X"00",
20151=>X"00",
20152=>X"00",
20153=>X"00",
20154=>X"00",
20155=>X"00",
20156=>X"00",
20157=>X"00",
20158=>X"00",
20159=>X"00",
20160=>X"00",
20161=>X"00",
20162=>X"00",
20163=>X"00",
20164=>X"00",
20165=>X"00",
20166=>X"00",
20167=>X"00",
20168=>X"00",
20169=>X"00",
20170=>X"00",
20171=>X"00",
20172=>X"00",
20173=>X"00",
20174=>X"00",
20175=>X"00",
20176=>X"00",
20177=>X"00",
20178=>X"00",
20179=>X"00",
20180=>X"00",
20181=>X"00",
20182=>X"00",
20183=>X"00",
20184=>X"00",
20185=>X"00",
20186=>X"00",
20187=>X"00",
20188=>X"00",
20189=>X"00",
20190=>X"00",
20191=>X"00",
20192=>X"00",
20193=>X"00",
20194=>X"00",
20195=>X"00",
20196=>X"00",
20197=>X"00",
20198=>X"00",
20199=>X"00",
20200=>X"00",
20201=>X"00",
20202=>X"00",
20203=>X"00",
20204=>X"00",
20205=>X"00",
20206=>X"00",
20207=>X"00",
20208=>X"00",
20209=>X"00",
20210=>X"00",
20211=>X"00",
20212=>X"00",
20213=>X"00",
20214=>X"00",
20215=>X"00",
20216=>X"00",
20217=>X"00",
20218=>X"00",
20219=>X"00",
20220=>X"00",
20221=>X"00",
20222=>X"00",
20223=>X"00",
20224=>X"00",
20225=>X"00",
20226=>X"00",
20227=>X"00",
20228=>X"00",
20229=>X"00",
20230=>X"00",
20231=>X"00",
20232=>X"00",
20233=>X"00",
20234=>X"00",
20235=>X"00",
20236=>X"00",
20237=>X"00",
20238=>X"00",
20239=>X"00",
20240=>X"00",
20241=>X"00",
20242=>X"00",
20243=>X"00",
20244=>X"00",
20245=>X"00",
20246=>X"00",
20247=>X"00",
20248=>X"00",
20249=>X"00",
20250=>X"00",
20251=>X"00",
20252=>X"00",
20253=>X"00",
20254=>X"00",
20255=>X"00",
20256=>X"00",
20257=>X"00",
20258=>X"00",
20259=>X"00",
20260=>X"00",
20261=>X"00",
20262=>X"00",
20263=>X"00",
20264=>X"00",
20265=>X"00",
20266=>X"00",
20267=>X"00",
20268=>X"00",
20269=>X"00",
20270=>X"00",
20271=>X"00",
20272=>X"00",
20273=>X"00",
20274=>X"00",
20275=>X"00",
20276=>X"00",
20277=>X"00",
20278=>X"00",
20279=>X"00",
20280=>X"00",
20281=>X"00",
20282=>X"00",
20283=>X"00",
20284=>X"00",
20285=>X"00",
20286=>X"00",
20287=>X"00",
20288=>X"00",
20289=>X"00",
20290=>X"00",
20291=>X"00",
20292=>X"00",
20293=>X"00",
20294=>X"00",
20295=>X"00",
20296=>X"00",
20297=>X"00",
20298=>X"00",
20299=>X"00",
20300=>X"00",
20301=>X"00",
20302=>X"00",
20303=>X"00",
20304=>X"00",
20305=>X"00",
20306=>X"00",
20307=>X"00",
20308=>X"00",
20309=>X"00",
20310=>X"00",
20311=>X"00",
20312=>X"00",
20313=>X"00",
20314=>X"00",
20315=>X"00",
20316=>X"00",
20317=>X"00",
20318=>X"00",
20319=>X"00",
20320=>X"00",
20321=>X"00",
20322=>X"00",
20323=>X"00",
20324=>X"00",
20325=>X"00",
20326=>X"00",
20327=>X"00",
20328=>X"00",
20329=>X"00",
20330=>X"00",
20331=>X"00",
20332=>X"00",
20333=>X"00",
20334=>X"00",
20335=>X"00",
20336=>X"00",
20337=>X"00",
20338=>X"00",
20339=>X"00",
20340=>X"00",
20341=>X"00",
20342=>X"00",
20343=>X"00",
20344=>X"00",
20345=>X"00",
20346=>X"00",
20347=>X"00",
20348=>X"00",
20349=>X"00",
20350=>X"00",
20351=>X"00",
20352=>X"00",
20353=>X"00",
20354=>X"00",
20355=>X"00",
20356=>X"00",
20357=>X"00",
20358=>X"00",
20359=>X"00",
20360=>X"00",
20361=>X"00",
20362=>X"00",
20363=>X"00",
20364=>X"00",
20365=>X"00",
20366=>X"00",
20367=>X"00",
20368=>X"00",
20369=>X"00",
20370=>X"00",
20371=>X"00",
20372=>X"00",
20373=>X"00",
20374=>X"00",
20375=>X"00",
20376=>X"00",
20377=>X"00",
20378=>X"00",
20379=>X"00",
20380=>X"00",
20381=>X"00",
20382=>X"00",
20383=>X"00",
20384=>X"00",
20385=>X"00",
20386=>X"00",
20387=>X"00",
20388=>X"00",
20389=>X"00",
20390=>X"00",
20391=>X"00",
20392=>X"00",
20393=>X"00",
20394=>X"00",
20395=>X"00",
20396=>X"00",
20397=>X"00",
20398=>X"00",
20399=>X"00",
20400=>X"00",
20401=>X"00",
20402=>X"00",
20403=>X"00",
20404=>X"00",
20405=>X"00",
20406=>X"00",
20407=>X"00",
20408=>X"00",
20409=>X"00",
20410=>X"00",
20411=>X"00",
20412=>X"00",
20413=>X"00",
20414=>X"00",
20415=>X"00",
20416=>X"00",
20417=>X"00",
20418=>X"00",
20419=>X"00",
20420=>X"00",
20421=>X"00",
20422=>X"00",
20423=>X"00",
20424=>X"00",
20425=>X"00",
20426=>X"00",
20427=>X"00",
20428=>X"00",
20429=>X"00",
20430=>X"00",
20431=>X"00",
20432=>X"00",
20433=>X"00",
20434=>X"00",
20435=>X"00",
20436=>X"00",
20437=>X"00",
20438=>X"00",
20439=>X"00",
20440=>X"00",
20441=>X"00",
20442=>X"00",
20443=>X"00",
20444=>X"00",
20445=>X"00",
20446=>X"00",
20447=>X"00",
20448=>X"00",
20449=>X"00",
20450=>X"00",
20451=>X"00",
20452=>X"00",
20453=>X"00",
20454=>X"00",
20455=>X"00",
20456=>X"00",
20457=>X"00",
20458=>X"00",
20459=>X"00",
20460=>X"00",
20461=>X"00",
20462=>X"00",
20463=>X"00",
20464=>X"00",
20465=>X"00",
20466=>X"00",
20467=>X"00",
20468=>X"00",
20469=>X"00",
20470=>X"00",
20471=>X"00",
20472=>X"00",
20473=>X"00",
20474=>X"00",
20475=>X"00",
20476=>X"00",
20477=>X"00",
20478=>X"00",
20479=>X"00",
20480=>X"00",
20481=>X"00",
20482=>X"00",
20483=>X"00",
20484=>X"00",
20485=>X"00",
20486=>X"00",
20487=>X"00",
20488=>X"00",
20489=>X"00",
20490=>X"00",
20491=>X"00",
20492=>X"00",
20493=>X"00",
20494=>X"00",
20495=>X"00",
20496=>X"00",
20497=>X"00",
20498=>X"00",
20499=>X"00",
20500=>X"00",
20501=>X"00",
20502=>X"00",
20503=>X"00",
20504=>X"00",
20505=>X"00",
20506=>X"00",
20507=>X"00",
20508=>X"00",
20509=>X"00",
20510=>X"00",
20511=>X"00",
20512=>X"00",
20513=>X"00",
20514=>X"00",
20515=>X"00",
20516=>X"00",
20517=>X"00",
20518=>X"00",
20519=>X"00",
20520=>X"00",
20521=>X"00",
20522=>X"00",
20523=>X"00",
20524=>X"00",
20525=>X"00",
20526=>X"00",
20527=>X"00",
20528=>X"00",
20529=>X"00",
20530=>X"00",
20531=>X"00",
20532=>X"00",
20533=>X"00",
20534=>X"00",
20535=>X"00",
20536=>X"00",
20537=>X"00",
20538=>X"00",
20539=>X"00",
20540=>X"00",
20541=>X"00",
20542=>X"00",
20543=>X"00",
20544=>X"00",
20545=>X"00",
20546=>X"00",
20547=>X"00",
20548=>X"00",
20549=>X"00",
20550=>X"00",
20551=>X"00",
20552=>X"00",
20553=>X"00",
20554=>X"00",
20555=>X"00",
20556=>X"00",
20557=>X"00",
20558=>X"00",
20559=>X"00",
20560=>X"00",
20561=>X"00",
20562=>X"00",
20563=>X"00",
20564=>X"00",
20565=>X"00",
20566=>X"00",
20567=>X"00",
20568=>X"00",
20569=>X"00",
20570=>X"00",
20571=>X"00",
20572=>X"00",
20573=>X"00",
20574=>X"00",
20575=>X"00",
20576=>X"00",
20577=>X"00",
20578=>X"00",
20579=>X"00",
20580=>X"00",
20581=>X"00",
20582=>X"00",
20583=>X"00",
20584=>X"00",
20585=>X"00",
20586=>X"00",
20587=>X"00",
20588=>X"00",
20589=>X"00",
20590=>X"00",
20591=>X"00",
20592=>X"00",
20593=>X"00",
20594=>X"00",
20595=>X"00",
20596=>X"00",
20597=>X"00",
20598=>X"00",
20599=>X"00",
20600=>X"00",
20601=>X"00",
20602=>X"00",
20603=>X"00",
20604=>X"00",
20605=>X"00",
20606=>X"00",
20607=>X"00",
20608=>X"00",
20609=>X"00",
20610=>X"00",
20611=>X"00",
20612=>X"00",
20613=>X"00",
20614=>X"00",
20615=>X"00",
20616=>X"00",
20617=>X"00",
20618=>X"00",
20619=>X"00",
20620=>X"00",
20621=>X"00",
20622=>X"00",
20623=>X"00",
20624=>X"00",
20625=>X"00",
20626=>X"00",
20627=>X"00",
20628=>X"00",
20629=>X"00",
20630=>X"00",
20631=>X"00",
20632=>X"00",
20633=>X"00",
20634=>X"00",
20635=>X"00",
20636=>X"00",
20637=>X"00",
20638=>X"00",
20639=>X"00",
20640=>X"00",
20641=>X"00",
20642=>X"00",
20643=>X"00",
20644=>X"00",
20645=>X"00",
20646=>X"00",
20647=>X"00",
20648=>X"00",
20649=>X"00",
20650=>X"00",
20651=>X"00",
20652=>X"00",
20653=>X"00",
20654=>X"00",
20655=>X"00",
20656=>X"00",
20657=>X"00",
20658=>X"00",
20659=>X"00",
20660=>X"00",
20661=>X"00",
20662=>X"00",
20663=>X"00",
20664=>X"00",
20665=>X"00",
20666=>X"00",
20667=>X"00",
20668=>X"00",
20669=>X"00",
20670=>X"00",
20671=>X"00",
20672=>X"00",
20673=>X"00",
20674=>X"00",
20675=>X"00",
20676=>X"00",
20677=>X"00",
20678=>X"00",
20679=>X"00",
20680=>X"00",
20681=>X"00",
20682=>X"00",
20683=>X"00",
20684=>X"00",
20685=>X"00",
20686=>X"00",
20687=>X"00",
20688=>X"00",
20689=>X"00",
20690=>X"00",
20691=>X"00",
20692=>X"00",
20693=>X"00",
20694=>X"00",
20695=>X"00",
20696=>X"00",
20697=>X"00",
20698=>X"00",
20699=>X"00",
20700=>X"00",
20701=>X"00",
20702=>X"00",
20703=>X"00",
20704=>X"00",
20705=>X"00",
20706=>X"00",
20707=>X"00",
20708=>X"00",
20709=>X"00",
20710=>X"00",
20711=>X"00",
20712=>X"00",
20713=>X"00",
20714=>X"00",
20715=>X"00",
20716=>X"00",
20717=>X"00",
20718=>X"00",
20719=>X"00",
20720=>X"00",
20721=>X"00",
20722=>X"00",
20723=>X"00",
20724=>X"00",
20725=>X"00",
20726=>X"00",
20727=>X"00",
20728=>X"00",
20729=>X"00",
20730=>X"00",
20731=>X"00",
20732=>X"00",
20733=>X"00",
20734=>X"00",
20735=>X"00",
20736=>X"00",
20737=>X"00",
20738=>X"00",
20739=>X"00",
20740=>X"00",
20741=>X"00",
20742=>X"00",
20743=>X"00",
20744=>X"00",
20745=>X"00",
20746=>X"00",
20747=>X"00",
20748=>X"00",
20749=>X"00",
20750=>X"00",
20751=>X"00",
20752=>X"00",
20753=>X"00",
20754=>X"00",
20755=>X"00",
20756=>X"00",
20757=>X"00",
20758=>X"00",
20759=>X"00",
20760=>X"00",
20761=>X"00",
20762=>X"00",
20763=>X"00",
20764=>X"00",
20765=>X"00",
20766=>X"00",
20767=>X"00",
20768=>X"00",
20769=>X"00",
20770=>X"00",
20771=>X"00",
20772=>X"00",
20773=>X"00",
20774=>X"00",
20775=>X"00",
20776=>X"00",
20777=>X"00",
20778=>X"00",
20779=>X"00",
20780=>X"00",
20781=>X"00",
20782=>X"00",
20783=>X"00",
20784=>X"00",
20785=>X"00",
20786=>X"00",
20787=>X"00",
20788=>X"00",
20789=>X"00",
20790=>X"00",
20791=>X"00",
20792=>X"00",
20793=>X"00",
20794=>X"00",
20795=>X"00",
20796=>X"00",
20797=>X"00",
20798=>X"00",
20799=>X"00",
20800=>X"00",
20801=>X"00",
20802=>X"00",
20803=>X"00",
20804=>X"00",
20805=>X"00",
20806=>X"00",
20807=>X"00",
20808=>X"00",
20809=>X"00",
20810=>X"00",
20811=>X"00",
20812=>X"00",
20813=>X"00",
20814=>X"00",
20815=>X"00",
20816=>X"00",
20817=>X"00",
20818=>X"00",
20819=>X"00",
20820=>X"00",
20821=>X"00",
20822=>X"00",
20823=>X"00",
20824=>X"00",
20825=>X"00",
20826=>X"00",
20827=>X"00",
20828=>X"00",
20829=>X"00",
20830=>X"00",
20831=>X"00",
20832=>X"00",
20833=>X"00",
20834=>X"00",
20835=>X"00",
20836=>X"00",
20837=>X"00",
20838=>X"00",
20839=>X"00",
20840=>X"00",
20841=>X"00",
20842=>X"00",
20843=>X"00",
20844=>X"00",
20845=>X"00",
20846=>X"00",
20847=>X"00",
20848=>X"00",
20849=>X"00",
20850=>X"00",
20851=>X"00",
20852=>X"00",
20853=>X"00",
20854=>X"00",
20855=>X"00",
20856=>X"00",
20857=>X"00",
20858=>X"00",
20859=>X"00",
20860=>X"00",
20861=>X"00",
20862=>X"00",
20863=>X"00",
20864=>X"00",
20865=>X"00",
20866=>X"00",
20867=>X"00",
20868=>X"00",
20869=>X"00",
20870=>X"00",
20871=>X"00",
20872=>X"00",
20873=>X"00",
20874=>X"00",
20875=>X"00",
20876=>X"00",
20877=>X"00",
20878=>X"00",
20879=>X"00",
20880=>X"00",
20881=>X"00",
20882=>X"00",
20883=>X"00",
20884=>X"00",
20885=>X"00",
20886=>X"00",
20887=>X"00",
20888=>X"00",
20889=>X"00",
20890=>X"00",
20891=>X"00",
20892=>X"00",
20893=>X"00",
20894=>X"00",
20895=>X"00",
20896=>X"00",
20897=>X"00",
20898=>X"00",
20899=>X"00",
20900=>X"00",
20901=>X"00",
20902=>X"00",
20903=>X"00",
20904=>X"00",
20905=>X"00",
20906=>X"00",
20907=>X"00",
20908=>X"00",
20909=>X"00",
20910=>X"00",
20911=>X"00",
20912=>X"00",
20913=>X"00",
20914=>X"00",
20915=>X"00",
20916=>X"00",
20917=>X"00",
20918=>X"00",
20919=>X"00",
20920=>X"00",
20921=>X"00",
20922=>X"00",
20923=>X"00",
20924=>X"00",
20925=>X"00",
20926=>X"00",
20927=>X"00",
20928=>X"00",
20929=>X"00",
20930=>X"00",
20931=>X"00",
20932=>X"00",
20933=>X"00",
20934=>X"00",
20935=>X"00",
20936=>X"00",
20937=>X"00",
20938=>X"00",
20939=>X"00",
20940=>X"00",
20941=>X"00",
20942=>X"00",
20943=>X"00",
20944=>X"00",
20945=>X"00",
20946=>X"00",
20947=>X"00",
20948=>X"00",
20949=>X"00",
20950=>X"00",
20951=>X"00",
20952=>X"00",
20953=>X"00",
20954=>X"00",
20955=>X"00",
20956=>X"00",
20957=>X"00",
20958=>X"00",
20959=>X"00",
20960=>X"00",
20961=>X"00",
20962=>X"00",
20963=>X"00",
20964=>X"00",
20965=>X"00",
20966=>X"00",
20967=>X"00",
20968=>X"00",
20969=>X"00",
20970=>X"00",
20971=>X"00",
20972=>X"00",
20973=>X"00",
20974=>X"00",
20975=>X"00",
20976=>X"00",
20977=>X"00",
20978=>X"00",
20979=>X"00",
20980=>X"00",
20981=>X"00",
20982=>X"00",
20983=>X"00",
20984=>X"00",
20985=>X"00",
20986=>X"00",
20987=>X"00",
20988=>X"00",
20989=>X"00",
20990=>X"00",
20991=>X"00",
20992=>X"00",
20993=>X"00",
20994=>X"00",
20995=>X"00",
20996=>X"00",
20997=>X"00",
20998=>X"00",
20999=>X"00",
21000=>X"00",
21001=>X"00",
21002=>X"00",
21003=>X"00",
21004=>X"00",
21005=>X"00",
21006=>X"00",
21007=>X"00",
21008=>X"00",
21009=>X"00",
21010=>X"00",
21011=>X"00",
21012=>X"00",
21013=>X"00",
21014=>X"00",
21015=>X"00",
21016=>X"00",
21017=>X"00",
21018=>X"00",
21019=>X"00",
21020=>X"00",
21021=>X"00",
21022=>X"00",
21023=>X"00",
21024=>X"00",
21025=>X"00",
21026=>X"00",
21027=>X"00",
21028=>X"00",
21029=>X"00",
21030=>X"00",
21031=>X"00",
21032=>X"00",
21033=>X"00",
21034=>X"00",
21035=>X"00",
21036=>X"00",
21037=>X"00",
21038=>X"00",
21039=>X"00",
21040=>X"00",
21041=>X"00",
21042=>X"00",
21043=>X"00",
21044=>X"00",
21045=>X"00",
21046=>X"00",
21047=>X"00",
21048=>X"00",
21049=>X"00",
21050=>X"00",
21051=>X"00",
21052=>X"00",
21053=>X"00",
21054=>X"00",
21055=>X"00",
21056=>X"00",
21057=>X"00",
21058=>X"00",
21059=>X"00",
21060=>X"00",
21061=>X"00",
21062=>X"00",
21063=>X"00",
21064=>X"00",
21065=>X"00",
21066=>X"00",
21067=>X"00",
21068=>X"00",
21069=>X"00",
21070=>X"00",
21071=>X"00",
21072=>X"00",
21073=>X"00",
21074=>X"00",
21075=>X"00",
21076=>X"00",
21077=>X"00",
21078=>X"00",
21079=>X"00",
21080=>X"00",
21081=>X"00",
21082=>X"00",
21083=>X"00",
21084=>X"00",
21085=>X"00",
21086=>X"00",
21087=>X"00",
21088=>X"00",
21089=>X"00",
21090=>X"00",
21091=>X"00",
21092=>X"00",
21093=>X"00",
21094=>X"00",
21095=>X"00",
21096=>X"00",
21097=>X"00",
21098=>X"00",
21099=>X"00",
21100=>X"00",
21101=>X"00",
21102=>X"00",
21103=>X"00",
21104=>X"00",
21105=>X"00",
21106=>X"00",
21107=>X"00",
21108=>X"00",
21109=>X"00",
21110=>X"00",
21111=>X"00",
21112=>X"00",
21113=>X"00",
21114=>X"00",
21115=>X"00",
21116=>X"00",
21117=>X"00",
21118=>X"00",
21119=>X"00",
21120=>X"00",
21121=>X"00",
21122=>X"00",
21123=>X"00",
21124=>X"00",
21125=>X"00",
21126=>X"00",
21127=>X"00",
21128=>X"00",
21129=>X"00",
21130=>X"00",
21131=>X"00",
21132=>X"00",
21133=>X"00",
21134=>X"00",
21135=>X"00",
21136=>X"00",
21137=>X"00",
21138=>X"00",
21139=>X"00",
21140=>X"00",
21141=>X"00",
21142=>X"00",
21143=>X"00",
21144=>X"00",
21145=>X"00",
21146=>X"00",
21147=>X"00",
21148=>X"00",
21149=>X"00",
21150=>X"00",
21151=>X"00",
21152=>X"00",
21153=>X"00",
21154=>X"00",
21155=>X"00",
21156=>X"00",
21157=>X"00",
21158=>X"00",
21159=>X"00",
21160=>X"00",
21161=>X"00",
21162=>X"00",
21163=>X"00",
21164=>X"00",
21165=>X"00",
21166=>X"00",
21167=>X"00",
21168=>X"00",
21169=>X"00",
21170=>X"00",
21171=>X"00",
21172=>X"00",
21173=>X"00",
21174=>X"00",
21175=>X"00",
21176=>X"00",
21177=>X"00",
21178=>X"00",
21179=>X"00",
21180=>X"00",
21181=>X"00",
21182=>X"00",
21183=>X"00",
21184=>X"00",
21185=>X"00",
21186=>X"00",
21187=>X"00",
21188=>X"00",
21189=>X"00",
21190=>X"00",
21191=>X"00",
21192=>X"00",
21193=>X"00",
21194=>X"00",
21195=>X"00",
21196=>X"00",
21197=>X"00",
21198=>X"00",
21199=>X"00",
21200=>X"00",
21201=>X"00",
21202=>X"00",
21203=>X"00",
21204=>X"00",
21205=>X"00",
21206=>X"00",
21207=>X"00",
21208=>X"00",
21209=>X"00",
21210=>X"00",
21211=>X"00",
21212=>X"00",
21213=>X"00",
21214=>X"00",
21215=>X"00",
21216=>X"00",
21217=>X"00",
21218=>X"00",
21219=>X"00",
21220=>X"00",
21221=>X"00",
21222=>X"00",
21223=>X"00",
21224=>X"00",
21225=>X"00",
21226=>X"00",
21227=>X"00",
21228=>X"00",
21229=>X"00",
21230=>X"00",
21231=>X"00",
21232=>X"00",
21233=>X"00",
21234=>X"00",
21235=>X"00",
21236=>X"00",
21237=>X"00",
21238=>X"00",
21239=>X"00",
21240=>X"00",
21241=>X"00",
21242=>X"00",
21243=>X"00",
21244=>X"00",
21245=>X"00",
21246=>X"00",
21247=>X"00",
21248=>X"00",
21249=>X"00",
21250=>X"00",
21251=>X"00",
21252=>X"00",
21253=>X"00",
21254=>X"00",
21255=>X"00",
21256=>X"00",
21257=>X"00",
21258=>X"00",
21259=>X"00",
21260=>X"00",
21261=>X"00",
21262=>X"00",
21263=>X"00",
21264=>X"00",
21265=>X"00",
21266=>X"00",
21267=>X"00",
21268=>X"00",
21269=>X"00",
21270=>X"00",
21271=>X"00",
21272=>X"00",
21273=>X"00",
21274=>X"00",
21275=>X"00",
21276=>X"00",
21277=>X"00",
21278=>X"00",
21279=>X"00",
21280=>X"00",
21281=>X"00",
21282=>X"00",
21283=>X"00",
21284=>X"00",
21285=>X"00",
21286=>X"00",
21287=>X"00",
21288=>X"00",
21289=>X"00",
21290=>X"00",
21291=>X"00",
21292=>X"00",
21293=>X"00",
21294=>X"00",
21295=>X"00",
21296=>X"00",
21297=>X"00",
21298=>X"00",
21299=>X"00",
21300=>X"00",
21301=>X"00",
21302=>X"00",
21303=>X"00",
21304=>X"00",
21305=>X"00",
21306=>X"00",
21307=>X"00",
21308=>X"00",
21309=>X"00",
21310=>X"00",
21311=>X"00",
21312=>X"00",
21313=>X"00",
21314=>X"00",
21315=>X"00",
21316=>X"00",
21317=>X"00",
21318=>X"00",
21319=>X"00",
21320=>X"00",
21321=>X"00",
21322=>X"00",
21323=>X"00",
21324=>X"00",
21325=>X"00",
21326=>X"00",
21327=>X"00",
21328=>X"00",
21329=>X"00",
21330=>X"00",
21331=>X"00",
21332=>X"00",
21333=>X"00",
21334=>X"00",
21335=>X"00",
21336=>X"00",
21337=>X"00",
21338=>X"00",
21339=>X"00",
21340=>X"00",
21341=>X"00",
21342=>X"00",
21343=>X"00",
21344=>X"00",
21345=>X"00",
21346=>X"00",
21347=>X"00",
21348=>X"00",
21349=>X"00",
21350=>X"00",
21351=>X"00",
21352=>X"00",
21353=>X"00",
21354=>X"00",
21355=>X"00",
21356=>X"00",
21357=>X"00",
21358=>X"00",
21359=>X"00",
21360=>X"00",
21361=>X"00",
21362=>X"00",
21363=>X"00",
21364=>X"00",
21365=>X"00",
21366=>X"00",
21367=>X"00",
21368=>X"00",
21369=>X"00",
21370=>X"00",
21371=>X"00",
21372=>X"00",
21373=>X"00",
21374=>X"00",
21375=>X"00",
21376=>X"00",
21377=>X"00",
21378=>X"00",
21379=>X"00",
21380=>X"00",
21381=>X"00",
21382=>X"00",
21383=>X"00",
21384=>X"00",
21385=>X"00",
21386=>X"00",
21387=>X"00",
21388=>X"00",
21389=>X"00",
21390=>X"00",
21391=>X"00",
21392=>X"00",
21393=>X"00",
21394=>X"00",
21395=>X"00",
21396=>X"00",
21397=>X"00",
21398=>X"00",
21399=>X"00",
21400=>X"00",
21401=>X"00",
21402=>X"00",
21403=>X"00",
21404=>X"00",
21405=>X"00",
21406=>X"00",
21407=>X"00",
21408=>X"00",
21409=>X"00",
21410=>X"00",
21411=>X"00",
21412=>X"00",
21413=>X"00",
21414=>X"00",
21415=>X"00",
21416=>X"00",
21417=>X"00",
21418=>X"00",
21419=>X"00",
21420=>X"00",
21421=>X"00",
21422=>X"00",
21423=>X"00",
21424=>X"00",
21425=>X"00",
21426=>X"00",
21427=>X"00",
21428=>X"00",
21429=>X"00",
21430=>X"00",
21431=>X"00",
21432=>X"00",
21433=>X"00",
21434=>X"00",
21435=>X"00",
21436=>X"00",
21437=>X"00",
21438=>X"00",
21439=>X"00",
21440=>X"00",
21441=>X"00",
21442=>X"00",
21443=>X"00",
21444=>X"00",
21445=>X"00",
21446=>X"00",
21447=>X"00",
21448=>X"00",
21449=>X"00",
21450=>X"00",
21451=>X"00",
21452=>X"00",
21453=>X"00",
21454=>X"00",
21455=>X"00",
21456=>X"00",
21457=>X"00",
21458=>X"00",
21459=>X"00",
21460=>X"00",
21461=>X"00",
21462=>X"00",
21463=>X"00",
21464=>X"00",
21465=>X"00",
21466=>X"00",
21467=>X"00",
21468=>X"00",
21469=>X"00",
21470=>X"00",
21471=>X"00",
21472=>X"00",
21473=>X"00",
21474=>X"00",
21475=>X"00",
21476=>X"00",
21477=>X"00",
21478=>X"00",
21479=>X"00",
21480=>X"00",
21481=>X"00",
21482=>X"00",
21483=>X"00",
21484=>X"00",
21485=>X"00",
21486=>X"00",
21487=>X"00",
21488=>X"00",
21489=>X"00",
21490=>X"00",
21491=>X"00",
21492=>X"00",
21493=>X"00",
21494=>X"00",
21495=>X"00",
21496=>X"00",
21497=>X"00",
21498=>X"00",
21499=>X"00",
21500=>X"00",
21501=>X"00",
21502=>X"00",
21503=>X"00",
21504=>X"00",
21505=>X"00",
21506=>X"00",
21507=>X"00",
21508=>X"00",
21509=>X"00",
21510=>X"00",
21511=>X"00",
21512=>X"00",
21513=>X"00",
21514=>X"00",
21515=>X"00",
21516=>X"00",
21517=>X"00",
21518=>X"00",
21519=>X"00",
21520=>X"00",
21521=>X"00",
21522=>X"00",
21523=>X"00",
21524=>X"00",
21525=>X"00",
21526=>X"00",
21527=>X"00",
21528=>X"00",
21529=>X"00",
21530=>X"00",
21531=>X"00",
21532=>X"00",
21533=>X"00",
21534=>X"00",
21535=>X"00",
21536=>X"00",
21537=>X"00",
21538=>X"00",
21539=>X"00",
21540=>X"00",
21541=>X"00",
21542=>X"00",
21543=>X"00",
21544=>X"00",
21545=>X"00",
21546=>X"00",
21547=>X"00",
21548=>X"00",
21549=>X"00",
21550=>X"00",
21551=>X"00",
21552=>X"00",
21553=>X"00",
21554=>X"00",
21555=>X"00",
21556=>X"00",
21557=>X"00",
21558=>X"00",
21559=>X"00",
21560=>X"00",
21561=>X"00",
21562=>X"00",
21563=>X"00",
21564=>X"00",
21565=>X"00",
21566=>X"00",
21567=>X"00",
21568=>X"00",
21569=>X"00",
21570=>X"00",
21571=>X"00",
21572=>X"00",
21573=>X"00",
21574=>X"00",
21575=>X"00",
21576=>X"00",
21577=>X"00",
21578=>X"00",
21579=>X"00",
21580=>X"00",
21581=>X"00",
21582=>X"00",
21583=>X"00",
21584=>X"00",
21585=>X"00",
21586=>X"00",
21587=>X"00",
21588=>X"00",
21589=>X"00",
21590=>X"00",
21591=>X"00",
21592=>X"00",
21593=>X"00",
21594=>X"00",
21595=>X"00",
21596=>X"00",
21597=>X"00",
21598=>X"00",
21599=>X"00",
21600=>X"00",
21601=>X"00",
21602=>X"00",
21603=>X"00",
21604=>X"00",
21605=>X"00",
21606=>X"00",
21607=>X"00",
21608=>X"00",
21609=>X"00",
21610=>X"00",
21611=>X"00",
21612=>X"00",
21613=>X"00",
21614=>X"00",
21615=>X"00",
21616=>X"00",
21617=>X"00",
21618=>X"00",
21619=>X"00",
21620=>X"00",
21621=>X"00",
21622=>X"00",
21623=>X"00",
21624=>X"00",
21625=>X"00",
21626=>X"00",
21627=>X"00",
21628=>X"00",
21629=>X"00",
21630=>X"00",
21631=>X"00",
21632=>X"00",
21633=>X"00",
21634=>X"00",
21635=>X"00",
21636=>X"00",
21637=>X"00",
21638=>X"00",
21639=>X"00",
21640=>X"00",
21641=>X"00",
21642=>X"00",
21643=>X"00",
21644=>X"00",
21645=>X"00",
21646=>X"00",
21647=>X"00",
21648=>X"00",
21649=>X"00",
21650=>X"00",
21651=>X"00",
21652=>X"00",
21653=>X"00",
21654=>X"00",
21655=>X"00",
21656=>X"00",
21657=>X"00",
21658=>X"00",
21659=>X"00",
21660=>X"00",
21661=>X"00",
21662=>X"00",
21663=>X"00",
21664=>X"00",
21665=>X"00",
21666=>X"00",
21667=>X"00",
21668=>X"00",
21669=>X"00",
21670=>X"00",
21671=>X"00",
21672=>X"00",
21673=>X"00",
21674=>X"00",
21675=>X"00",
21676=>X"00",
21677=>X"00",
21678=>X"00",
21679=>X"00",
21680=>X"00",
21681=>X"00",
21682=>X"00",
21683=>X"00",
21684=>X"00",
21685=>X"00",
21686=>X"00",
21687=>X"00",
21688=>X"00",
21689=>X"00",
21690=>X"00",
21691=>X"00",
21692=>X"00",
21693=>X"00",
21694=>X"00",
21695=>X"00",
21696=>X"00",
21697=>X"00",
21698=>X"00",
21699=>X"00",
21700=>X"00",
21701=>X"00",
21702=>X"00",
21703=>X"00",
21704=>X"00",
21705=>X"00",
21706=>X"00",
21707=>X"00",
21708=>X"00",
21709=>X"00",
21710=>X"00",
21711=>X"00",
21712=>X"00",
21713=>X"00",
21714=>X"00",
21715=>X"00",
21716=>X"00",
21717=>X"00",
21718=>X"00",
21719=>X"00",
21720=>X"00",
21721=>X"00",
21722=>X"00",
21723=>X"00",
21724=>X"00",
21725=>X"00",
21726=>X"00",
21727=>X"00",
21728=>X"00",
21729=>X"00",
21730=>X"00",
21731=>X"00",
21732=>X"00",
21733=>X"00",
21734=>X"00",
21735=>X"00",
21736=>X"00",
21737=>X"00",
21738=>X"00",
21739=>X"00",
21740=>X"00",
21741=>X"00",
21742=>X"00",
21743=>X"00",
21744=>X"00",
21745=>X"00",
21746=>X"00",
21747=>X"00",
21748=>X"00",
21749=>X"00",
21750=>X"00",
21751=>X"00",
21752=>X"00",
21753=>X"00",
21754=>X"00",
21755=>X"00",
21756=>X"00",
21757=>X"00",
21758=>X"00",
21759=>X"00",
21760=>X"00",
21761=>X"00",
21762=>X"00",
21763=>X"00",
21764=>X"00",
21765=>X"00",
21766=>X"00",
21767=>X"00",
21768=>X"00",
21769=>X"00",
21770=>X"00",
21771=>X"00",
21772=>X"00",
21773=>X"00",
21774=>X"00",
21775=>X"00",
21776=>X"00",
21777=>X"00",
21778=>X"00",
21779=>X"00",
21780=>X"00",
21781=>X"00",
21782=>X"00",
21783=>X"00",
21784=>X"00",
21785=>X"00",
21786=>X"00",
21787=>X"00",
21788=>X"00",
21789=>X"00",
21790=>X"00",
21791=>X"00",
21792=>X"00",
21793=>X"00",
21794=>X"00",
21795=>X"00",
21796=>X"00",
21797=>X"00",
21798=>X"00",
21799=>X"00",
21800=>X"00",
21801=>X"00",
21802=>X"00",
21803=>X"00",
21804=>X"00",
21805=>X"00",
21806=>X"00",
21807=>X"00",
21808=>X"00",
21809=>X"00",
21810=>X"00",
21811=>X"00",
21812=>X"00",
21813=>X"00",
21814=>X"00",
21815=>X"00",
21816=>X"00",
21817=>X"00",
21818=>X"00",
21819=>X"00",
21820=>X"00",
21821=>X"00",
21822=>X"00",
21823=>X"00",
21824=>X"00",
21825=>X"00",
21826=>X"00",
21827=>X"00",
21828=>X"00",
21829=>X"00",
21830=>X"00",
21831=>X"00",
21832=>X"00",
21833=>X"00",
21834=>X"00",
21835=>X"00",
21836=>X"00",
21837=>X"00",
21838=>X"00",
21839=>X"00",
21840=>X"00",
21841=>X"00",
21842=>X"00",
21843=>X"00",
21844=>X"00",
21845=>X"00",
21846=>X"00",
21847=>X"00",
21848=>X"00",
21849=>X"00",
21850=>X"00",
21851=>X"00",
21852=>X"00",
21853=>X"00",
21854=>X"00",
21855=>X"00",
21856=>X"00",
21857=>X"00",
21858=>X"00",
21859=>X"00",
21860=>X"00",
21861=>X"00",
21862=>X"00",
21863=>X"00",
21864=>X"00",
21865=>X"00",
21866=>X"00",
21867=>X"00",
21868=>X"00",
21869=>X"00",
21870=>X"00",
21871=>X"00",
21872=>X"00",
21873=>X"00",
21874=>X"00",
21875=>X"00",
21876=>X"00",
21877=>X"00",
21878=>X"00",
21879=>X"00",
21880=>X"00",
21881=>X"00",
21882=>X"00",
21883=>X"00",
21884=>X"00",
21885=>X"00",
21886=>X"00",
21887=>X"00",
21888=>X"00",
21889=>X"00",
21890=>X"00",
21891=>X"00",
21892=>X"00",
21893=>X"00",
21894=>X"00",
21895=>X"00",
21896=>X"00",
21897=>X"00",
21898=>X"00",
21899=>X"00",
21900=>X"00",
21901=>X"00",
21902=>X"00",
21903=>X"00",
21904=>X"00",
21905=>X"00",
21906=>X"00",
21907=>X"00",
21908=>X"00",
21909=>X"00",
21910=>X"00",
21911=>X"00",
21912=>X"00",
21913=>X"00",
21914=>X"00",
21915=>X"00",
21916=>X"00",
21917=>X"00",
21918=>X"00",
21919=>X"00",
21920=>X"00",
21921=>X"00",
21922=>X"00",
21923=>X"00",
21924=>X"00",
21925=>X"00",
21926=>X"00",
21927=>X"00",
21928=>X"00",
21929=>X"00",
21930=>X"00",
21931=>X"00",
21932=>X"00",
21933=>X"00",
21934=>X"00",
21935=>X"00",
21936=>X"00",
21937=>X"00",
21938=>X"00",
21939=>X"00",
21940=>X"00",
21941=>X"00",
21942=>X"00",
21943=>X"00",
21944=>X"00",
21945=>X"00",
21946=>X"00",
21947=>X"00",
21948=>X"00",
21949=>X"00",
21950=>X"00",
21951=>X"00",
21952=>X"00",
21953=>X"00",
21954=>X"00",
21955=>X"00",
21956=>X"00",
21957=>X"00",
21958=>X"00",
21959=>X"00",
21960=>X"00",
21961=>X"00",
21962=>X"00",
21963=>X"00",
21964=>X"00",
21965=>X"00",
21966=>X"00",
21967=>X"00",
21968=>X"00",
21969=>X"00",
21970=>X"00",
21971=>X"00",
21972=>X"00",
21973=>X"00",
21974=>X"00",
21975=>X"00",
21976=>X"00",
21977=>X"00",
21978=>X"00",
21979=>X"00",
21980=>X"00",
21981=>X"00",
21982=>X"00",
21983=>X"00",
21984=>X"00",
21985=>X"00",
21986=>X"00",
21987=>X"00",
21988=>X"00",
21989=>X"00",
21990=>X"00",
21991=>X"00",
21992=>X"00",
21993=>X"00",
21994=>X"00",
21995=>X"00",
21996=>X"00",
21997=>X"00",
21998=>X"00",
21999=>X"00",
22000=>X"00",
22001=>X"00",
22002=>X"00",
22003=>X"00",
22004=>X"00",
22005=>X"00",
22006=>X"00",
22007=>X"00",
22008=>X"00",
22009=>X"00",
22010=>X"00",
22011=>X"00",
22012=>X"00",
22013=>X"00",
22014=>X"00",
22015=>X"00",
22016=>X"00",
22017=>X"00",
22018=>X"00",
22019=>X"00",
22020=>X"00",
22021=>X"00",
22022=>X"00",
22023=>X"00",
22024=>X"00",
22025=>X"00",
22026=>X"00",
22027=>X"00",
22028=>X"00",
22029=>X"00",
22030=>X"00",
22031=>X"00",
22032=>X"00",
22033=>X"00",
22034=>X"00",
22035=>X"00",
22036=>X"00",
22037=>X"00",
22038=>X"00",
22039=>X"00",
22040=>X"00",
22041=>X"00",
22042=>X"00",
22043=>X"00",
22044=>X"00",
22045=>X"00",
22046=>X"00",
22047=>X"00",
22048=>X"00",
22049=>X"00",
22050=>X"00",
22051=>X"00",
22052=>X"00",
22053=>X"00",
22054=>X"00",
22055=>X"00",
22056=>X"00",
22057=>X"00",
22058=>X"00",
22059=>X"00",
22060=>X"00",
22061=>X"00",
22062=>X"00",
22063=>X"00",
22064=>X"00",
22065=>X"00",
22066=>X"00",
22067=>X"00",
22068=>X"00",
22069=>X"00",
22070=>X"00",
22071=>X"00",
22072=>X"00",
22073=>X"00",
22074=>X"00",
22075=>X"00",
22076=>X"00",
22077=>X"00",
22078=>X"00",
22079=>X"00",
22080=>X"00",
22081=>X"00",
22082=>X"00",
22083=>X"00",
22084=>X"00",
22085=>X"00",
22086=>X"00",
22087=>X"00",
22088=>X"00",
22089=>X"00",
22090=>X"00",
22091=>X"00",
22092=>X"00",
22093=>X"00",
22094=>X"00",
22095=>X"00",
22096=>X"00",
22097=>X"00",
22098=>X"00",
22099=>X"00",
22100=>X"00",
22101=>X"00",
22102=>X"00",
22103=>X"00",
22104=>X"00",
22105=>X"00",
22106=>X"00",
22107=>X"00",
22108=>X"00",
22109=>X"00",
22110=>X"00",
22111=>X"00",
22112=>X"00",
22113=>X"00",
22114=>X"00",
22115=>X"00",
22116=>X"00",
22117=>X"00",
22118=>X"00",
22119=>X"00",
22120=>X"00",
22121=>X"00",
22122=>X"00",
22123=>X"00",
22124=>X"00",
22125=>X"00",
22126=>X"00",
22127=>X"00",
22128=>X"00",
22129=>X"00",
22130=>X"00",
22131=>X"00",
22132=>X"00",
22133=>X"00",
22134=>X"00",
22135=>X"00",
22136=>X"00",
22137=>X"00",
22138=>X"00",
22139=>X"00",
22140=>X"00",
22141=>X"00",
22142=>X"00",
22143=>X"00",
22144=>X"00",
22145=>X"00",
22146=>X"00",
22147=>X"00",
22148=>X"00",
22149=>X"00",
22150=>X"00",
22151=>X"00",
22152=>X"00",
22153=>X"00",
22154=>X"00",
22155=>X"00",
22156=>X"00",
22157=>X"00",
22158=>X"00",
22159=>X"00",
22160=>X"00",
22161=>X"00",
22162=>X"00",
22163=>X"00",
22164=>X"00",
22165=>X"00",
22166=>X"00",
22167=>X"00",
22168=>X"00",
22169=>X"00",
22170=>X"00",
22171=>X"00",
22172=>X"00",
22173=>X"00",
22174=>X"00",
22175=>X"00",
22176=>X"00",
22177=>X"00",
22178=>X"00",
22179=>X"00",
22180=>X"00",
22181=>X"00",
22182=>X"00",
22183=>X"00",
22184=>X"00",
22185=>X"00",
22186=>X"00",
22187=>X"00",
22188=>X"00",
22189=>X"00",
22190=>X"00",
22191=>X"00",
22192=>X"00",
22193=>X"00",
22194=>X"00",
22195=>X"00",
22196=>X"00",
22197=>X"00",
22198=>X"00",
22199=>X"00",
22200=>X"00",
22201=>X"00",
22202=>X"00",
22203=>X"00",
22204=>X"00",
22205=>X"00",
22206=>X"00",
22207=>X"00",
22208=>X"00",
22209=>X"00",
22210=>X"00",
22211=>X"00",
22212=>X"00",
22213=>X"00",
22214=>X"00",
22215=>X"00",
22216=>X"00",
22217=>X"00",
22218=>X"00",
22219=>X"00",
22220=>X"00",
22221=>X"00",
22222=>X"00",
22223=>X"00",
22224=>X"00",
22225=>X"00",
22226=>X"00",
22227=>X"00",
22228=>X"00",
22229=>X"00",
22230=>X"00",
22231=>X"00",
22232=>X"00",
22233=>X"00",
22234=>X"00",
22235=>X"00",
22236=>X"00",
22237=>X"00",
22238=>X"00",
22239=>X"00",
22240=>X"00",
22241=>X"00",
22242=>X"00",
22243=>X"00",
22244=>X"00",
22245=>X"00",
22246=>X"00",
22247=>X"00",
22248=>X"00",
22249=>X"00",
22250=>X"00",
22251=>X"00",
22252=>X"00",
22253=>X"00",
22254=>X"00",
22255=>X"00",
22256=>X"00",
22257=>X"00",
22258=>X"00",
22259=>X"00",
22260=>X"00",
22261=>X"00",
22262=>X"00",
22263=>X"00",
22264=>X"00",
22265=>X"00",
22266=>X"00",
22267=>X"00",
22268=>X"00",
22269=>X"00",
22270=>X"00",
22271=>X"00",
22272=>X"00",
22273=>X"00",
22274=>X"00",
22275=>X"00",
22276=>X"00",
22277=>X"00",
22278=>X"00",
22279=>X"00",
22280=>X"00",
22281=>X"00",
22282=>X"00",
22283=>X"00",
22284=>X"00",
22285=>X"00",
22286=>X"00",
22287=>X"00",
22288=>X"00",
22289=>X"00",
22290=>X"00",
22291=>X"00",
22292=>X"00",
22293=>X"00",
22294=>X"00",
22295=>X"00",
22296=>X"00",
22297=>X"00",
22298=>X"00",
22299=>X"00",
22300=>X"00",
22301=>X"00",
22302=>X"00",
22303=>X"00",
22304=>X"00",
22305=>X"00",
22306=>X"00",
22307=>X"00",
22308=>X"00",
22309=>X"00",
22310=>X"00",
22311=>X"00",
22312=>X"00",
22313=>X"00",
22314=>X"00",
22315=>X"00",
22316=>X"00",
22317=>X"00",
22318=>X"00",
22319=>X"00",
22320=>X"00",
22321=>X"00",
22322=>X"00",
22323=>X"00",
22324=>X"00",
22325=>X"00",
22326=>X"00",
22327=>X"00",
22328=>X"00",
22329=>X"00",
22330=>X"00",
22331=>X"00",
22332=>X"00",
22333=>X"00",
22334=>X"00",
22335=>X"00",
22336=>X"00",
22337=>X"00",
22338=>X"00",
22339=>X"00",
22340=>X"00",
22341=>X"00",
22342=>X"00",
22343=>X"00",
22344=>X"00",
22345=>X"00",
22346=>X"00",
22347=>X"00",
22348=>X"00",
22349=>X"00",
22350=>X"00",
22351=>X"00",
22352=>X"00",
22353=>X"00",
22354=>X"00",
22355=>X"00",
22356=>X"00",
22357=>X"00",
22358=>X"00",
22359=>X"00",
22360=>X"00",
22361=>X"00",
22362=>X"00",
22363=>X"00",
22364=>X"00",
22365=>X"00",
22366=>X"00",
22367=>X"00",
22368=>X"00",
22369=>X"00",
22370=>X"00",
22371=>X"00",
22372=>X"00",
22373=>X"00",
22374=>X"00",
22375=>X"00",
22376=>X"00",
22377=>X"00",
22378=>X"00",
22379=>X"00",
22380=>X"00",
22381=>X"00",
22382=>X"00",
22383=>X"00",
22384=>X"00",
22385=>X"00",
22386=>X"00",
22387=>X"00",
22388=>X"00",
22389=>X"00",
22390=>X"00",
22391=>X"00",
22392=>X"00",
22393=>X"00",
22394=>X"00",
22395=>X"00",
22396=>X"00",
22397=>X"00",
22398=>X"00",
22399=>X"00",
22400=>X"00",
22401=>X"00",
22402=>X"00",
22403=>X"00",
22404=>X"00",
22405=>X"00",
22406=>X"00",
22407=>X"00",
22408=>X"00",
22409=>X"00",
22410=>X"00",
22411=>X"00",
22412=>X"00",
22413=>X"00",
22414=>X"00",
22415=>X"00",
22416=>X"00",
22417=>X"00",
22418=>X"00",
22419=>X"00",
22420=>X"00",
22421=>X"00",
22422=>X"00",
22423=>X"00",
22424=>X"00",
22425=>X"00",
22426=>X"00",
22427=>X"00",
22428=>X"00",
22429=>X"00",
22430=>X"00",
22431=>X"00",
22432=>X"00",
22433=>X"00",
22434=>X"00",
22435=>X"00",
22436=>X"00",
22437=>X"00",
22438=>X"00",
22439=>X"00",
22440=>X"00",
22441=>X"00",
22442=>X"00",
22443=>X"00",
22444=>X"00",
22445=>X"00",
22446=>X"00",
22447=>X"00",
22448=>X"00",
22449=>X"00",
22450=>X"00",
22451=>X"00",
22452=>X"00",
22453=>X"00",
22454=>X"00",
22455=>X"00",
22456=>X"00",
22457=>X"00",
22458=>X"00",
22459=>X"00",
22460=>X"00",
22461=>X"00",
22462=>X"00",
22463=>X"00",
22464=>X"00",
22465=>X"00",
22466=>X"00",
22467=>X"00",
22468=>X"00",
22469=>X"00",
22470=>X"00",
22471=>X"00",
22472=>X"00",
22473=>X"00",
22474=>X"00",
22475=>X"00",
22476=>X"00",
22477=>X"00",
22478=>X"00",
22479=>X"00",
22480=>X"00",
22481=>X"00",
22482=>X"00",
22483=>X"00",
22484=>X"00",
22485=>X"00",
22486=>X"00",
22487=>X"00",
22488=>X"00",
22489=>X"00",
22490=>X"00",
22491=>X"00",
22492=>X"00",
22493=>X"00",
22494=>X"00",
22495=>X"00",
22496=>X"00",
22497=>X"00",
22498=>X"00",
22499=>X"00",
22500=>X"00",
22501=>X"00",
22502=>X"00",
22503=>X"00",
22504=>X"00",
22505=>X"00",
22506=>X"00",
22507=>X"00",
22508=>X"00",
22509=>X"00",
22510=>X"00",
22511=>X"00",
22512=>X"00",
22513=>X"00",
22514=>X"00",
22515=>X"00",
22516=>X"00",
22517=>X"00",
22518=>X"00",
22519=>X"00",
22520=>X"00",
22521=>X"00",
22522=>X"00",
22523=>X"00",
22524=>X"00",
22525=>X"00",
22526=>X"00",
22527=>X"00",
22528=>X"00",
22529=>X"00",
22530=>X"00",
22531=>X"00",
22532=>X"00",
22533=>X"00",
22534=>X"00",
22535=>X"00",
22536=>X"00",
22537=>X"00",
22538=>X"00",
22539=>X"00",
22540=>X"00",
22541=>X"00",
22542=>X"00",
22543=>X"00",
22544=>X"00",
22545=>X"00",
22546=>X"00",
22547=>X"00",
22548=>X"00",
22549=>X"00",
22550=>X"00",
22551=>X"00",
22552=>X"00",
22553=>X"00",
22554=>X"00",
22555=>X"00",
22556=>X"00",
22557=>X"00",
22558=>X"00",
22559=>X"00",
22560=>X"00",
22561=>X"00",
22562=>X"00",
22563=>X"00",
22564=>X"00",
22565=>X"00",
22566=>X"00",
22567=>X"00",
22568=>X"00",
22569=>X"00",
22570=>X"00",
22571=>X"00",
22572=>X"00",
22573=>X"00",
22574=>X"00",
22575=>X"00",
22576=>X"00",
22577=>X"00",
22578=>X"00",
22579=>X"00",
22580=>X"00",
22581=>X"00",
22582=>X"00",
22583=>X"00",
22584=>X"00",
22585=>X"00",
22586=>X"00",
22587=>X"00",
22588=>X"00",
22589=>X"00",
22590=>X"00",
22591=>X"00",
22592=>X"00",
22593=>X"00",
22594=>X"00",
22595=>X"00",
22596=>X"00",
22597=>X"00",
22598=>X"00",
22599=>X"00",
22600=>X"00",
22601=>X"00",
22602=>X"00",
22603=>X"00",
22604=>X"00",
22605=>X"00",
22606=>X"00",
22607=>X"00",
22608=>X"00",
22609=>X"00",
22610=>X"00",
22611=>X"00",
22612=>X"00",
22613=>X"00",
22614=>X"00",
22615=>X"00",
22616=>X"00",
22617=>X"00",
22618=>X"00",
22619=>X"00",
22620=>X"00",
22621=>X"00",
22622=>X"00",
22623=>X"00",
22624=>X"00",
22625=>X"00",
22626=>X"00",
22627=>X"00",
22628=>X"00",
22629=>X"00",
22630=>X"00",
22631=>X"00",
22632=>X"00",
22633=>X"00",
22634=>X"00",
22635=>X"00",
22636=>X"00",
22637=>X"00",
22638=>X"00",
22639=>X"00",
22640=>X"00",
22641=>X"00",
22642=>X"00",
22643=>X"00",
22644=>X"00",
22645=>X"00",
22646=>X"00",
22647=>X"00",
22648=>X"00",
22649=>X"00",
22650=>X"00",
22651=>X"00",
22652=>X"00",
22653=>X"00",
22654=>X"00",
22655=>X"00",
22656=>X"00",
22657=>X"00",
22658=>X"00",
22659=>X"00",
22660=>X"00",
22661=>X"00",
22662=>X"00",
22663=>X"00",
22664=>X"00",
22665=>X"00",
22666=>X"00",
22667=>X"00",
22668=>X"00",
22669=>X"00",
22670=>X"00",
22671=>X"00",
22672=>X"00",
22673=>X"00",
22674=>X"00",
22675=>X"00",
22676=>X"00",
22677=>X"00",
22678=>X"00",
22679=>X"00",
22680=>X"00",
22681=>X"00",
22682=>X"00",
22683=>X"00",
22684=>X"00",
22685=>X"00",
22686=>X"00",
22687=>X"00",
22688=>X"00",
22689=>X"00",
22690=>X"00",
22691=>X"00",
22692=>X"00",
22693=>X"00",
22694=>X"00",
22695=>X"00",
22696=>X"00",
22697=>X"00",
22698=>X"00",
22699=>X"00",
22700=>X"00",
22701=>X"00",
22702=>X"00",
22703=>X"00",
22704=>X"00",
22705=>X"00",
22706=>X"00",
22707=>X"00",
22708=>X"00",
22709=>X"00",
22710=>X"00",
22711=>X"00",
22712=>X"00",
22713=>X"00",
22714=>X"00",
22715=>X"00",
22716=>X"00",
22717=>X"00",
22718=>X"00",
22719=>X"00",
22720=>X"00",
22721=>X"00",
22722=>X"00",
22723=>X"00",
22724=>X"00",
22725=>X"00",
22726=>X"00",
22727=>X"00",
22728=>X"00",
22729=>X"00",
22730=>X"00",
22731=>X"00",
22732=>X"00",
22733=>X"00",
22734=>X"00",
22735=>X"00",
22736=>X"00",
22737=>X"00",
22738=>X"00",
22739=>X"00",
22740=>X"00",
22741=>X"00",
22742=>X"00",
22743=>X"00",
22744=>X"00",
22745=>X"00",
22746=>X"00",
22747=>X"00",
22748=>X"00",
22749=>X"00",
22750=>X"00",
22751=>X"00",
22752=>X"00",
22753=>X"00",
22754=>X"00",
22755=>X"00",
22756=>X"00",
22757=>X"00",
22758=>X"00",
22759=>X"00",
22760=>X"00",
22761=>X"00",
22762=>X"00",
22763=>X"00",
22764=>X"00",
22765=>X"00",
22766=>X"00",
22767=>X"00",
22768=>X"00",
22769=>X"00",
22770=>X"00",
22771=>X"00",
22772=>X"00",
22773=>X"00",
22774=>X"00",
22775=>X"00",
22776=>X"00",
22777=>X"00",
22778=>X"00",
22779=>X"00",
22780=>X"00",
22781=>X"00",
22782=>X"00",
22783=>X"00",
22784=>X"00",
22785=>X"00",
22786=>X"00",
22787=>X"00",
22788=>X"00",
22789=>X"00",
22790=>X"00",
22791=>X"00",
22792=>X"00",
22793=>X"00",
22794=>X"00",
22795=>X"00",
22796=>X"00",
22797=>X"00",
22798=>X"00",
22799=>X"00",
22800=>X"00",
22801=>X"00",
22802=>X"00",
22803=>X"00",
22804=>X"00",
22805=>X"00",
22806=>X"00",
22807=>X"00",
22808=>X"00",
22809=>X"00",
22810=>X"00",
22811=>X"00",
22812=>X"00",
22813=>X"00",
22814=>X"00",
22815=>X"00",
22816=>X"00",
22817=>X"00",
22818=>X"00",
22819=>X"00",
22820=>X"00",
22821=>X"00",
22822=>X"00",
22823=>X"00",
22824=>X"00",
22825=>X"00",
22826=>X"00",
22827=>X"00",
22828=>X"00",
22829=>X"00",
22830=>X"00",
22831=>X"00",
22832=>X"00",
22833=>X"00",
22834=>X"00",
22835=>X"00",
22836=>X"00",
22837=>X"00",
22838=>X"00",
22839=>X"00",
22840=>X"00",
22841=>X"00",
22842=>X"00",
22843=>X"00",
22844=>X"00",
22845=>X"00",
22846=>X"00",
22847=>X"00",
22848=>X"00",
22849=>X"00",
22850=>X"00",
22851=>X"00",
22852=>X"00",
22853=>X"00",
22854=>X"00",
22855=>X"00",
22856=>X"00",
22857=>X"00",
22858=>X"00",
22859=>X"00",
22860=>X"00",
22861=>X"00",
22862=>X"00",
22863=>X"00",
22864=>X"00",
22865=>X"00",
22866=>X"00",
22867=>X"00",
22868=>X"00",
22869=>X"00",
22870=>X"00",
22871=>X"00",
22872=>X"00",
22873=>X"00",
22874=>X"00",
22875=>X"00",
22876=>X"00",
22877=>X"00",
22878=>X"00",
22879=>X"00",
22880=>X"00",
22881=>X"00",
22882=>X"00",
22883=>X"00",
22884=>X"00",
22885=>X"00",
22886=>X"00",
22887=>X"00",
22888=>X"00",
22889=>X"00",
22890=>X"00",
22891=>X"00",
22892=>X"00",
22893=>X"00",
22894=>X"00",
22895=>X"00",
22896=>X"00",
22897=>X"00",
22898=>X"00",
22899=>X"00",
22900=>X"00",
22901=>X"00",
22902=>X"00",
22903=>X"00",
22904=>X"00",
22905=>X"00",
22906=>X"00",
22907=>X"00",
22908=>X"00",
22909=>X"00",
22910=>X"00",
22911=>X"00",
22912=>X"00",
22913=>X"00",
22914=>X"00",
22915=>X"00",
22916=>X"00",
22917=>X"00",
22918=>X"00",
22919=>X"00",
22920=>X"00",
22921=>X"00",
22922=>X"00",
22923=>X"00",
22924=>X"00",
22925=>X"00",
22926=>X"00",
22927=>X"00",
22928=>X"00",
22929=>X"00",
22930=>X"00",
22931=>X"00",
22932=>X"00",
22933=>X"00",
22934=>X"00",
22935=>X"00",
22936=>X"00",
22937=>X"00",
22938=>X"00",
22939=>X"00",
22940=>X"00",
22941=>X"00",
22942=>X"00",
22943=>X"00",
22944=>X"00",
22945=>X"00",
22946=>X"00",
22947=>X"00",
22948=>X"00",
22949=>X"00",
22950=>X"00",
22951=>X"00",
22952=>X"00",
22953=>X"00",
22954=>X"00",
22955=>X"00",
22956=>X"00",
22957=>X"00",
22958=>X"00",
22959=>X"00",
22960=>X"00",
22961=>X"00",
22962=>X"00",
22963=>X"00",
22964=>X"00",
22965=>X"00",
22966=>X"00",
22967=>X"00",
22968=>X"00",
22969=>X"00",
22970=>X"00",
22971=>X"00",
22972=>X"00",
22973=>X"00",
22974=>X"00",
22975=>X"00",
22976=>X"00",
22977=>X"00",
22978=>X"00",
22979=>X"00",
22980=>X"00",
22981=>X"00",
22982=>X"00",
22983=>X"00",
22984=>X"00",
22985=>X"00",
22986=>X"00",
22987=>X"00",
22988=>X"00",
22989=>X"00",
22990=>X"00",
22991=>X"00",
22992=>X"00",
22993=>X"00",
22994=>X"00",
22995=>X"00",
22996=>X"00",
22997=>X"00",
22998=>X"00",
22999=>X"00",
23000=>X"00",
23001=>X"00",
23002=>X"00",
23003=>X"00",
23004=>X"00",
23005=>X"00",
23006=>X"00",
23007=>X"00",
23008=>X"00",
23009=>X"00",
23010=>X"00",
23011=>X"00",
23012=>X"00",
23013=>X"00",
23014=>X"00",
23015=>X"00",
23016=>X"00",
23017=>X"00",
23018=>X"00",
23019=>X"00",
23020=>X"00",
23021=>X"00",
23022=>X"00",
23023=>X"00",
23024=>X"00",
23025=>X"00",
23026=>X"00",
23027=>X"00",
23028=>X"00",
23029=>X"00",
23030=>X"00",
23031=>X"00",
23032=>X"00",
23033=>X"00",
23034=>X"00",
23035=>X"00",
23036=>X"00",
23037=>X"00",
23038=>X"00",
23039=>X"00",
23040=>X"00",
23041=>X"00",
23042=>X"00",
23043=>X"00",
23044=>X"00",
23045=>X"00",
23046=>X"00",
23047=>X"00",
23048=>X"00",
23049=>X"00",
23050=>X"00",
23051=>X"00",
23052=>X"00",
23053=>X"00",
23054=>X"00",
23055=>X"00",
23056=>X"00",
23057=>X"00",
23058=>X"00",
23059=>X"00",
23060=>X"00",
23061=>X"00",
23062=>X"00",
23063=>X"00",
23064=>X"00",
23065=>X"00",
23066=>X"00",
23067=>X"00",
23068=>X"00",
23069=>X"00",
23070=>X"00",
23071=>X"00",
23072=>X"00",
23073=>X"00",
23074=>X"00",
23075=>X"00",
23076=>X"00",
23077=>X"00",
23078=>X"00",
23079=>X"00",
23080=>X"00",
23081=>X"00",
23082=>X"00",
23083=>X"00",
23084=>X"00",
23085=>X"00",
23086=>X"00",
23087=>X"00",
23088=>X"00",
23089=>X"00",
23090=>X"00",
23091=>X"00",
23092=>X"00",
23093=>X"00",
23094=>X"00",
23095=>X"00",
23096=>X"00",
23097=>X"00",
23098=>X"00",
23099=>X"00",
23100=>X"00",
23101=>X"00",
23102=>X"00",
23103=>X"00",
23104=>X"00",
23105=>X"00",
23106=>X"00",
23107=>X"00",
23108=>X"00",
23109=>X"00",
23110=>X"00",
23111=>X"00",
23112=>X"00",
23113=>X"00",
23114=>X"00",
23115=>X"00",
23116=>X"00",
23117=>X"00",
23118=>X"00",
23119=>X"00",
23120=>X"00",
23121=>X"00",
23122=>X"00",
23123=>X"00",
23124=>X"00",
23125=>X"00",
23126=>X"00",
23127=>X"00",
23128=>X"00",
23129=>X"00",
23130=>X"00",
23131=>X"00",
23132=>X"00",
23133=>X"00",
23134=>X"00",
23135=>X"00",
23136=>X"00",
23137=>X"00",
23138=>X"00",
23139=>X"00",
23140=>X"00",
23141=>X"00",
23142=>X"00",
23143=>X"00",
23144=>X"00",
23145=>X"00",
23146=>X"00",
23147=>X"00",
23148=>X"00",
23149=>X"00",
23150=>X"00",
23151=>X"00",
23152=>X"00",
23153=>X"00",
23154=>X"00",
23155=>X"00",
23156=>X"00",
23157=>X"00",
23158=>X"00",
23159=>X"00",
23160=>X"00",
23161=>X"00",
23162=>X"00",
23163=>X"00",
23164=>X"00",
23165=>X"00",
23166=>X"00",
23167=>X"00",
23168=>X"00",
23169=>X"00",
23170=>X"00",
23171=>X"00",
23172=>X"00",
23173=>X"00",
23174=>X"00",
23175=>X"00",
23176=>X"00",
23177=>X"00",
23178=>X"00",
23179=>X"00",
23180=>X"00",
23181=>X"00",
23182=>X"00",
23183=>X"00",
23184=>X"00",
23185=>X"00",
23186=>X"00",
23187=>X"00",
23188=>X"00",
23189=>X"00",
23190=>X"00",
23191=>X"00",
23192=>X"00",
23193=>X"00",
23194=>X"00",
23195=>X"00",
23196=>X"00",
23197=>X"00",
23198=>X"00",
23199=>X"00",
23200=>X"00",
23201=>X"00",
23202=>X"00",
23203=>X"00",
23204=>X"00",
23205=>X"00",
23206=>X"00",
23207=>X"00",
23208=>X"00",
23209=>X"00",
23210=>X"00",
23211=>X"00",
23212=>X"00",
23213=>X"00",
23214=>X"00",
23215=>X"00",
23216=>X"00",
23217=>X"00",
23218=>X"00",
23219=>X"00",
23220=>X"00",
23221=>X"00",
23222=>X"00",
23223=>X"00",
23224=>X"00",
23225=>X"00",
23226=>X"00",
23227=>X"00",
23228=>X"00",
23229=>X"00",
23230=>X"00",
23231=>X"00",
23232=>X"00",
23233=>X"00",
23234=>X"00",
23235=>X"00",
23236=>X"00",
23237=>X"00",
23238=>X"00",
23239=>X"00",
23240=>X"00",
23241=>X"00",
23242=>X"00",
23243=>X"00",
23244=>X"00",
23245=>X"00",
23246=>X"00",
23247=>X"00",
23248=>X"00",
23249=>X"00",
23250=>X"00",
23251=>X"00",
23252=>X"00",
23253=>X"00",
23254=>X"00",
23255=>X"00",
23256=>X"00",
23257=>X"00",
23258=>X"00",
23259=>X"00",
23260=>X"00",
23261=>X"00",
23262=>X"00",
23263=>X"00",
23264=>X"00",
23265=>X"00",
23266=>X"00",
23267=>X"00",
23268=>X"00",
23269=>X"00",
23270=>X"00",
23271=>X"00",
23272=>X"00",
23273=>X"00",
23274=>X"00",
23275=>X"00",
23276=>X"00",
23277=>X"00",
23278=>X"00",
23279=>X"00",
23280=>X"00",
23281=>X"00",
23282=>X"00",
23283=>X"00",
23284=>X"00",
23285=>X"00",
23286=>X"00",
23287=>X"00",
23288=>X"00",
23289=>X"00",
23290=>X"00",
23291=>X"00",
23292=>X"00",
23293=>X"00",
23294=>X"00",
23295=>X"00",
23296=>X"00",
23297=>X"00",
23298=>X"00",
23299=>X"00",
23300=>X"00",
23301=>X"00",
23302=>X"00",
23303=>X"00",
23304=>X"00",
23305=>X"00",
23306=>X"00",
23307=>X"00",
23308=>X"00",
23309=>X"00",
23310=>X"00",
23311=>X"00",
23312=>X"00",
23313=>X"00",
23314=>X"00",
23315=>X"00",
23316=>X"00",
23317=>X"00",
23318=>X"00",
23319=>X"00",
23320=>X"00",
23321=>X"00",
23322=>X"00",
23323=>X"00",
23324=>X"00",
23325=>X"00",
23326=>X"00",
23327=>X"00",
23328=>X"00",
23329=>X"00",
23330=>X"00",
23331=>X"00",
23332=>X"00",
23333=>X"00",
23334=>X"00",
23335=>X"00",
23336=>X"00",
23337=>X"00",
23338=>X"00",
23339=>X"00",
23340=>X"00",
23341=>X"00",
23342=>X"00",
23343=>X"00",
23344=>X"00",
23345=>X"00",
23346=>X"00",
23347=>X"00",
23348=>X"00",
23349=>X"00",
23350=>X"00",
23351=>X"00",
23352=>X"00",
23353=>X"00",
23354=>X"00",
23355=>X"00",
23356=>X"00",
23357=>X"00",
23358=>X"00",
23359=>X"00",
23360=>X"00",
23361=>X"00",
23362=>X"00",
23363=>X"00",
23364=>X"00",
23365=>X"00",
23366=>X"00",
23367=>X"00",
23368=>X"00",
23369=>X"00",
23370=>X"00",
23371=>X"00",
23372=>X"00",
23373=>X"00",
23374=>X"00",
23375=>X"00",
23376=>X"00",
23377=>X"00",
23378=>X"00",
23379=>X"00",
23380=>X"00",
23381=>X"00",
23382=>X"00",
23383=>X"00",
23384=>X"00",
23385=>X"00",
23386=>X"00",
23387=>X"00",
23388=>X"00",
23389=>X"00",
23390=>X"00",
23391=>X"00",
23392=>X"00",
23393=>X"00",
23394=>X"00",
23395=>X"00",
23396=>X"00",
23397=>X"00",
23398=>X"00",
23399=>X"00",
23400=>X"00",
23401=>X"00",
23402=>X"00",
23403=>X"00",
23404=>X"00",
23405=>X"00",
23406=>X"00",
23407=>X"00",
23408=>X"00",
23409=>X"00",
23410=>X"00",
23411=>X"00",
23412=>X"00",
23413=>X"00",
23414=>X"00",
23415=>X"00",
23416=>X"00",
23417=>X"00",
23418=>X"00",
23419=>X"00",
23420=>X"00",
23421=>X"00",
23422=>X"00",
23423=>X"00",
23424=>X"00",
23425=>X"00",
23426=>X"00",
23427=>X"00",
23428=>X"00",
23429=>X"00",
23430=>X"00",
23431=>X"00",
23432=>X"00",
23433=>X"00",
23434=>X"00",
23435=>X"00",
23436=>X"00",
23437=>X"00",
23438=>X"00",
23439=>X"00",
23440=>X"00",
23441=>X"00",
23442=>X"00",
23443=>X"00",
23444=>X"00",
23445=>X"00",
23446=>X"00",
23447=>X"00",
23448=>X"00",
23449=>X"00",
23450=>X"00",
23451=>X"00",
23452=>X"00",
23453=>X"00",
23454=>X"00",
23455=>X"00",
23456=>X"00",
23457=>X"00",
23458=>X"00",
23459=>X"00",
23460=>X"00",
23461=>X"00",
23462=>X"00",
23463=>X"00",
23464=>X"00",
23465=>X"00",
23466=>X"00",
23467=>X"00",
23468=>X"00",
23469=>X"00",
23470=>X"00",
23471=>X"00",
23472=>X"00",
23473=>X"00",
23474=>X"00",
23475=>X"00",
23476=>X"00",
23477=>X"00",
23478=>X"00",
23479=>X"00",
23480=>X"00",
23481=>X"00",
23482=>X"00",
23483=>X"00",
23484=>X"00",
23485=>X"00",
23486=>X"00",
23487=>X"00",
23488=>X"00",
23489=>X"00",
23490=>X"00",
23491=>X"00",
23492=>X"00",
23493=>X"00",
23494=>X"00",
23495=>X"00",
23496=>X"00",
23497=>X"00",
23498=>X"00",
23499=>X"00",
23500=>X"00",
23501=>X"00",
23502=>X"00",
23503=>X"00",
23504=>X"00",
23505=>X"00",
23506=>X"00",
23507=>X"00",
23508=>X"00",
23509=>X"00",
23510=>X"00",
23511=>X"00",
23512=>X"00",
23513=>X"00",
23514=>X"00",
23515=>X"00",
23516=>X"00",
23517=>X"00",
23518=>X"00",
23519=>X"00",
23520=>X"00",
23521=>X"00",
23522=>X"00",
23523=>X"00",
23524=>X"00",
23525=>X"00",
23526=>X"00",
23527=>X"00",
23528=>X"00",
23529=>X"00",
23530=>X"00",
23531=>X"00",
23532=>X"00",
23533=>X"00",
23534=>X"00",
23535=>X"00",
23536=>X"00",
23537=>X"00",
23538=>X"00",
23539=>X"00",
23540=>X"00",
23541=>X"00",
23542=>X"00",
23543=>X"00",
23544=>X"00",
23545=>X"00",
23546=>X"00",
23547=>X"00",
23548=>X"00",
23549=>X"00",
23550=>X"00",
23551=>X"00",
23552=>X"00",
23553=>X"00",
23554=>X"00",
23555=>X"00",
23556=>X"00",
23557=>X"00",
23558=>X"00",
23559=>X"00",
23560=>X"00",
23561=>X"00",
23562=>X"00",
23563=>X"00",
23564=>X"00",
23565=>X"00",
23566=>X"00",
23567=>X"00",
23568=>X"00",
23569=>X"00",
23570=>X"00",
23571=>X"00",
23572=>X"00",
23573=>X"00",
23574=>X"00",
23575=>X"00",
23576=>X"00",
23577=>X"00",
23578=>X"00",
23579=>X"00",
23580=>X"00",
23581=>X"00",
23582=>X"00",
23583=>X"00",
23584=>X"00",
23585=>X"00",
23586=>X"00",
23587=>X"00",
23588=>X"00",
23589=>X"00",
23590=>X"00",
23591=>X"00",
23592=>X"00",
23593=>X"00",
23594=>X"00",
23595=>X"00",
23596=>X"00",
23597=>X"00",
23598=>X"00",
23599=>X"00",
23600=>X"00",
23601=>X"00",
23602=>X"00",
23603=>X"00",
23604=>X"00",
23605=>X"00",
23606=>X"00",
23607=>X"00",
23608=>X"00",
23609=>X"00",
23610=>X"00",
23611=>X"00",
23612=>X"00",
23613=>X"00",
23614=>X"00",
23615=>X"00",
23616=>X"00",
23617=>X"00",
23618=>X"00",
23619=>X"00",
23620=>X"00",
23621=>X"00",
23622=>X"00",
23623=>X"00",
23624=>X"00",
23625=>X"00",
23626=>X"00",
23627=>X"00",
23628=>X"00",
23629=>X"00",
23630=>X"00",
23631=>X"00",
23632=>X"00",
23633=>X"00",
23634=>X"00",
23635=>X"00",
23636=>X"00",
23637=>X"00",
23638=>X"00",
23639=>X"00",
23640=>X"00",
23641=>X"00",
23642=>X"00",
23643=>X"00",
23644=>X"00",
23645=>X"00",
23646=>X"00",
23647=>X"00",
23648=>X"00",
23649=>X"00",
23650=>X"00",
23651=>X"00",
23652=>X"00",
23653=>X"00",
23654=>X"00",
23655=>X"00",
23656=>X"00",
23657=>X"00",
23658=>X"00",
23659=>X"00",
23660=>X"00",
23661=>X"00",
23662=>X"00",
23663=>X"00",
23664=>X"00",
23665=>X"00",
23666=>X"00",
23667=>X"00",
23668=>X"00",
23669=>X"00",
23670=>X"00",
23671=>X"00",
23672=>X"00",
23673=>X"00",
23674=>X"00",
23675=>X"00",
23676=>X"00",
23677=>X"00",
23678=>X"00",
23679=>X"00",
23680=>X"00",
23681=>X"00",
23682=>X"00",
23683=>X"00",
23684=>X"00",
23685=>X"00",
23686=>X"00",
23687=>X"00",
23688=>X"00",
23689=>X"00",
23690=>X"00",
23691=>X"00",
23692=>X"00",
23693=>X"00",
23694=>X"00",
23695=>X"00",
23696=>X"00",
23697=>X"00",
23698=>X"00",
23699=>X"00",
23700=>X"00",
23701=>X"00",
23702=>X"00",
23703=>X"00",
23704=>X"00",
23705=>X"00",
23706=>X"00",
23707=>X"00",
23708=>X"00",
23709=>X"00",
23710=>X"00",
23711=>X"00",
23712=>X"00",
23713=>X"00",
23714=>X"00",
23715=>X"00",
23716=>X"00",
23717=>X"00",
23718=>X"00",
23719=>X"00",
23720=>X"00",
23721=>X"00",
23722=>X"00",
23723=>X"00",
23724=>X"00",
23725=>X"00",
23726=>X"00",
23727=>X"00",
23728=>X"00",
23729=>X"00",
23730=>X"00",
23731=>X"00",
23732=>X"00",
23733=>X"00",
23734=>X"00",
23735=>X"00",
23736=>X"00",
23737=>X"00",
23738=>X"00",
23739=>X"00",
23740=>X"00",
23741=>X"00",
23742=>X"00",
23743=>X"00",
23744=>X"00",
23745=>X"00",
23746=>X"00",
23747=>X"00",
23748=>X"00",
23749=>X"00",
23750=>X"00",
23751=>X"00",
23752=>X"00",
23753=>X"00",
23754=>X"00",
23755=>X"00",
23756=>X"00",
23757=>X"00",
23758=>X"00",
23759=>X"00",
23760=>X"00",
23761=>X"00",
23762=>X"00",
23763=>X"00",
23764=>X"00",
23765=>X"00",
23766=>X"00",
23767=>X"00",
23768=>X"00",
23769=>X"00",
23770=>X"00",
23771=>X"00",
23772=>X"00",
23773=>X"00",
23774=>X"00",
23775=>X"00",
23776=>X"00",
23777=>X"00",
23778=>X"00",
23779=>X"00",
23780=>X"00",
23781=>X"00",
23782=>X"00",
23783=>X"00",
23784=>X"00",
23785=>X"00",
23786=>X"00",
23787=>X"00",
23788=>X"00",
23789=>X"00",
23790=>X"00",
23791=>X"00",
23792=>X"00",
23793=>X"00",
23794=>X"00",
23795=>X"00",
23796=>X"00",
23797=>X"00",
23798=>X"00",
23799=>X"00",
23800=>X"00",
23801=>X"00",
23802=>X"00",
23803=>X"00",
23804=>X"00",
23805=>X"00",
23806=>X"00",
23807=>X"00",
23808=>X"00",
23809=>X"00",
23810=>X"00",
23811=>X"00",
23812=>X"00",
23813=>X"00",
23814=>X"00",
23815=>X"00",
23816=>X"00",
23817=>X"00",
23818=>X"00",
23819=>X"00",
23820=>X"00",
23821=>X"00",
23822=>X"00",
23823=>X"00",
23824=>X"00",
23825=>X"00",
23826=>X"00",
23827=>X"00",
23828=>X"00",
23829=>X"00",
23830=>X"00",
23831=>X"00",
23832=>X"00",
23833=>X"00",
23834=>X"00",
23835=>X"00",
23836=>X"00",
23837=>X"00",
23838=>X"00",
23839=>X"00",
23840=>X"00",
23841=>X"00",
23842=>X"00",
23843=>X"00",
23844=>X"00",
23845=>X"00",
23846=>X"00",
23847=>X"00",
23848=>X"00",
23849=>X"00",
23850=>X"00",
23851=>X"00",
23852=>X"00",
23853=>X"00",
23854=>X"00",
23855=>X"00",
23856=>X"00",
23857=>X"00",
23858=>X"00",
23859=>X"00",
23860=>X"00",
23861=>X"00",
23862=>X"00",
23863=>X"00",
23864=>X"00",
23865=>X"00",
23866=>X"00",
23867=>X"00",
23868=>X"00",
23869=>X"00",
23870=>X"00",
23871=>X"00",
23872=>X"00",
23873=>X"00",
23874=>X"00",
23875=>X"00",
23876=>X"00",
23877=>X"00",
23878=>X"00",
23879=>X"00",
23880=>X"00",
23881=>X"00",
23882=>X"00",
23883=>X"00",
23884=>X"00",
23885=>X"00",
23886=>X"00",
23887=>X"00",
23888=>X"00",
23889=>X"00",
23890=>X"00",
23891=>X"00",
23892=>X"00",
23893=>X"00",
23894=>X"00",
23895=>X"00",
23896=>X"00",
23897=>X"00",
23898=>X"00",
23899=>X"00",
23900=>X"00",
23901=>X"00",
23902=>X"00",
23903=>X"00",
23904=>X"00",
23905=>X"00",
23906=>X"00",
23907=>X"00",
23908=>X"00",
23909=>X"00",
23910=>X"00",
23911=>X"00",
23912=>X"00",
23913=>X"00",
23914=>X"00",
23915=>X"00",
23916=>X"00",
23917=>X"00",
23918=>X"00",
23919=>X"00",
23920=>X"00",
23921=>X"00",
23922=>X"00",
23923=>X"00",
23924=>X"00",
23925=>X"00",
23926=>X"00",
23927=>X"00",
23928=>X"00",
23929=>X"00",
23930=>X"00",
23931=>X"00",
23932=>X"00",
23933=>X"00",
23934=>X"00",
23935=>X"00",
23936=>X"00",
23937=>X"00",
23938=>X"00",
23939=>X"00",
23940=>X"00",
23941=>X"00",
23942=>X"00",
23943=>X"00",
23944=>X"00",
23945=>X"00",
23946=>X"00",
23947=>X"00",
23948=>X"00",
23949=>X"00",
23950=>X"00",
23951=>X"00",
23952=>X"00",
23953=>X"00",
23954=>X"00",
23955=>X"00",
23956=>X"00",
23957=>X"00",
23958=>X"00",
23959=>X"00",
23960=>X"00",
23961=>X"00",
23962=>X"00",
23963=>X"00",
23964=>X"00",
23965=>X"00",
23966=>X"00",
23967=>X"00",
23968=>X"00",
23969=>X"00",
23970=>X"00",
23971=>X"00",
23972=>X"00",
23973=>X"00",
23974=>X"00",
23975=>X"00",
23976=>X"00",
23977=>X"00",
23978=>X"00",
23979=>X"00",
23980=>X"00",
23981=>X"00",
23982=>X"00",
23983=>X"00",
23984=>X"00",
23985=>X"00",
23986=>X"00",
23987=>X"00",
23988=>X"00",
23989=>X"00",
23990=>X"00",
23991=>X"00",
23992=>X"00",
23993=>X"00",
23994=>X"00",
23995=>X"00",
23996=>X"00",
23997=>X"00",
23998=>X"00",
23999=>X"00",
24000=>X"00",
24001=>X"00",
24002=>X"00",
24003=>X"00",
24004=>X"00",
24005=>X"00",
24006=>X"00",
24007=>X"00",
24008=>X"00",
24009=>X"00",
24010=>X"00",
24011=>X"00",
24012=>X"00",
24013=>X"00",
24014=>X"00",
24015=>X"00",
24016=>X"00",
24017=>X"00",
24018=>X"00",
24019=>X"00",
24020=>X"00",
24021=>X"00",
24022=>X"00",
24023=>X"00",
24024=>X"00",
24025=>X"00",
24026=>X"00",
24027=>X"00",
24028=>X"00",
24029=>X"00",
24030=>X"00",
24031=>X"00",
24032=>X"00",
24033=>X"00",
24034=>X"00",
24035=>X"00",
24036=>X"00",
24037=>X"00",
24038=>X"00",
24039=>X"00",
24040=>X"00",
24041=>X"00",
24042=>X"00",
24043=>X"00",
24044=>X"00",
24045=>X"00",
24046=>X"00",
24047=>X"00",
24048=>X"00",
24049=>X"00",
24050=>X"00",
24051=>X"00",
24052=>X"00",
24053=>X"00",
24054=>X"00",
24055=>X"00",
24056=>X"00",
24057=>X"00",
24058=>X"00",
24059=>X"00",
24060=>X"00",
24061=>X"00",
24062=>X"00",
24063=>X"00",
24064=>X"00",
24065=>X"00",
24066=>X"00",
24067=>X"00",
24068=>X"00",
24069=>X"00",
24070=>X"00",
24071=>X"00",
24072=>X"00",
24073=>X"00",
24074=>X"00",
24075=>X"00",
24076=>X"00",
24077=>X"00",
24078=>X"00",
24079=>X"00",
24080=>X"00",
24081=>X"00",
24082=>X"00",
24083=>X"00",
24084=>X"00",
24085=>X"00",
24086=>X"00",
24087=>X"00",
24088=>X"00",
24089=>X"00",
24090=>X"00",
24091=>X"00",
24092=>X"00",
24093=>X"00",
24094=>X"00",
24095=>X"00",
24096=>X"00",
24097=>X"00",
24098=>X"00",
24099=>X"00",
24100=>X"00",
24101=>X"00",
24102=>X"00",
24103=>X"00",
24104=>X"00",
24105=>X"00",
24106=>X"00",
24107=>X"00",
24108=>X"00",
24109=>X"00",
24110=>X"00",
24111=>X"00",
24112=>X"00",
24113=>X"00",
24114=>X"00",
24115=>X"00",
24116=>X"00",
24117=>X"00",
24118=>X"00",
24119=>X"00",
24120=>X"00",
24121=>X"00",
24122=>X"00",
24123=>X"00",
24124=>X"00",
24125=>X"00",
24126=>X"00",
24127=>X"00",
24128=>X"00",
24129=>X"00",
24130=>X"00",
24131=>X"00",
24132=>X"00",
24133=>X"00",
24134=>X"00",
24135=>X"00",
24136=>X"00",
24137=>X"00",
24138=>X"00",
24139=>X"00",
24140=>X"00",
24141=>X"00",
24142=>X"00",
24143=>X"00",
24144=>X"00",
24145=>X"00",
24146=>X"00",
24147=>X"00",
24148=>X"00",
24149=>X"00",
24150=>X"00",
24151=>X"00",
24152=>X"00",
24153=>X"00",
24154=>X"00",
24155=>X"00",
24156=>X"00",
24157=>X"00",
24158=>X"00",
24159=>X"00",
24160=>X"00",
24161=>X"00",
24162=>X"00",
24163=>X"00",
24164=>X"00",
24165=>X"00",
24166=>X"00",
24167=>X"00",
24168=>X"00",
24169=>X"00",
24170=>X"00",
24171=>X"00",
24172=>X"00",
24173=>X"00",
24174=>X"00",
24175=>X"00",
24176=>X"00",
24177=>X"00",
24178=>X"00",
24179=>X"00",
24180=>X"00",
24181=>X"00",
24182=>X"00",
24183=>X"00",
24184=>X"00",
24185=>X"00",
24186=>X"00",
24187=>X"00",
24188=>X"00",
24189=>X"00",
24190=>X"00",
24191=>X"00",
24192=>X"00",
24193=>X"00",
24194=>X"00",
24195=>X"00",
24196=>X"00",
24197=>X"00",
24198=>X"00",
24199=>X"00",
24200=>X"00",
24201=>X"00",
24202=>X"00",
24203=>X"00",
24204=>X"00",
24205=>X"00",
24206=>X"00",
24207=>X"00",
24208=>X"00",
24209=>X"00",
24210=>X"00",
24211=>X"00",
24212=>X"00",
24213=>X"00",
24214=>X"00",
24215=>X"00",
24216=>X"00",
24217=>X"00",
24218=>X"00",
24219=>X"00",
24220=>X"00",
24221=>X"00",
24222=>X"00",
24223=>X"00",
24224=>X"00",
24225=>X"00",
24226=>X"00",
24227=>X"00",
24228=>X"00",
24229=>X"00",
24230=>X"00",
24231=>X"00",
24232=>X"00",
24233=>X"00",
24234=>X"00",
24235=>X"00",
24236=>X"00",
24237=>X"00",
24238=>X"00",
24239=>X"00",
24240=>X"00",
24241=>X"00",
24242=>X"00",
24243=>X"00",
24244=>X"00",
24245=>X"00",
24246=>X"00",
24247=>X"00",
24248=>X"00",
24249=>X"00",
24250=>X"00",
24251=>X"00",
24252=>X"00",
24253=>X"00",
24254=>X"00",
24255=>X"00",
24256=>X"00",
24257=>X"00",
24258=>X"00",
24259=>X"00",
24260=>X"00",
24261=>X"00",
24262=>X"00",
24263=>X"00",
24264=>X"00",
24265=>X"00",
24266=>X"00",
24267=>X"00",
24268=>X"00",
24269=>X"00",
24270=>X"00",
24271=>X"00",
24272=>X"00",
24273=>X"00",
24274=>X"00",
24275=>X"00",
24276=>X"00",
24277=>X"00",
24278=>X"00",
24279=>X"00",
24280=>X"00",
24281=>X"00",
24282=>X"00",
24283=>X"00",
24284=>X"00",
24285=>X"00",
24286=>X"00",
24287=>X"00",
24288=>X"00",
24289=>X"00",
24290=>X"00",
24291=>X"00",
24292=>X"00",
24293=>X"00",
24294=>X"00",
24295=>X"00",
24296=>X"00",
24297=>X"00",
24298=>X"00",
24299=>X"00",
24300=>X"00",
24301=>X"00",
24302=>X"00",
24303=>X"00",
24304=>X"00",
24305=>X"00",
24306=>X"00",
24307=>X"00",
24308=>X"00",
24309=>X"00",
24310=>X"00",
24311=>X"00",
24312=>X"00",
24313=>X"00",
24314=>X"00",
24315=>X"00",
24316=>X"00",
24317=>X"00",
24318=>X"00",
24319=>X"00",
24320=>X"00",
24321=>X"00",
24322=>X"00",
24323=>X"00",
24324=>X"00",
24325=>X"00",
24326=>X"00",
24327=>X"00",
24328=>X"00",
24329=>X"00",
24330=>X"00",
24331=>X"00",
24332=>X"00",
24333=>X"00",
24334=>X"00",
24335=>X"00",
24336=>X"00",
24337=>X"00",
24338=>X"00",
24339=>X"00",
24340=>X"00",
24341=>X"00",
24342=>X"00",
24343=>X"00",
24344=>X"00",
24345=>X"00",
24346=>X"00",
24347=>X"00",
24348=>X"00",
24349=>X"00",
24350=>X"00",
24351=>X"00",
24352=>X"00",
24353=>X"00",
24354=>X"00",
24355=>X"00",
24356=>X"00",
24357=>X"00",
24358=>X"00",
24359=>X"00",
24360=>X"00",
24361=>X"00",
24362=>X"00",
24363=>X"00",
24364=>X"00",
24365=>X"00",
24366=>X"00",
24367=>X"00",
24368=>X"00",
24369=>X"00",
24370=>X"00",
24371=>X"00",
24372=>X"00",
24373=>X"00",
24374=>X"00",
24375=>X"00",
24376=>X"00",
24377=>X"00",
24378=>X"00",
24379=>X"00",
24380=>X"00",
24381=>X"00",
24382=>X"00",
24383=>X"00",
24384=>X"00",
24385=>X"00",
24386=>X"00",
24387=>X"00",
24388=>X"00",
24389=>X"00",
24390=>X"00",
24391=>X"00",
24392=>X"00",
24393=>X"00",
24394=>X"00",
24395=>X"00",
24396=>X"00",
24397=>X"00",
24398=>X"00",
24399=>X"00",
24400=>X"00",
24401=>X"00",
24402=>X"00",
24403=>X"00",
24404=>X"00",
24405=>X"00",
24406=>X"00",
24407=>X"00",
24408=>X"00",
24409=>X"00",
24410=>X"00",
24411=>X"00",
24412=>X"00",
24413=>X"00",
24414=>X"00",
24415=>X"00",
24416=>X"00",
24417=>X"00",
24418=>X"00",
24419=>X"00",
24420=>X"00",
24421=>X"00",
24422=>X"00",
24423=>X"00",
24424=>X"00",
24425=>X"00",
24426=>X"00",
24427=>X"00",
24428=>X"00",
24429=>X"00",
24430=>X"00",
24431=>X"00",
24432=>X"00",
24433=>X"00",
24434=>X"00",
24435=>X"00",
24436=>X"00",
24437=>X"00",
24438=>X"00",
24439=>X"00",
24440=>X"00",
24441=>X"00",
24442=>X"00",
24443=>X"00",
24444=>X"00",
24445=>X"00",
24446=>X"00",
24447=>X"00",
24448=>X"00",
24449=>X"00",
24450=>X"00",
24451=>X"00",
24452=>X"00",
24453=>X"00",
24454=>X"00",
24455=>X"00",
24456=>X"00",
24457=>X"00",
24458=>X"00",
24459=>X"00",
24460=>X"00",
24461=>X"00",
24462=>X"00",
24463=>X"00",
24464=>X"00",
24465=>X"00",
24466=>X"00",
24467=>X"00",
24468=>X"00",
24469=>X"00",
24470=>X"00",
24471=>X"00",
24472=>X"00",
24473=>X"00",
24474=>X"00",
24475=>X"00",
24476=>X"00",
24477=>X"00",
24478=>X"00",
24479=>X"00",
24480=>X"00",
24481=>X"00",
24482=>X"00",
24483=>X"00",
24484=>X"00",
24485=>X"00",
24486=>X"00",
24487=>X"00",
24488=>X"00",
24489=>X"00",
24490=>X"00",
24491=>X"00",
24492=>X"00",
24493=>X"00",
24494=>X"00",
24495=>X"00",
24496=>X"00",
24497=>X"00",
24498=>X"00",
24499=>X"00",
24500=>X"00",
24501=>X"00",
24502=>X"00",
24503=>X"00",
24504=>X"00",
24505=>X"00",
24506=>X"00",
24507=>X"00",
24508=>X"00",
24509=>X"00",
24510=>X"00",
24511=>X"00",
24512=>X"00",
24513=>X"00",
24514=>X"00",
24515=>X"00",
24516=>X"00",
24517=>X"00",
24518=>X"00",
24519=>X"00",
24520=>X"00",
24521=>X"00",
24522=>X"00",
24523=>X"00",
24524=>X"00",
24525=>X"00",
24526=>X"00",
24527=>X"00",
24528=>X"00",
24529=>X"00",
24530=>X"00",
24531=>X"00",
24532=>X"00",
24533=>X"00",
24534=>X"00",
24535=>X"00",
24536=>X"00",
24537=>X"00",
24538=>X"00",
24539=>X"00",
24540=>X"00",
24541=>X"00",
24542=>X"00",
24543=>X"00",
24544=>X"00",
24545=>X"00",
24546=>X"00",
24547=>X"00",
24548=>X"00",
24549=>X"00",
24550=>X"00",
24551=>X"00",
24552=>X"00",
24553=>X"00",
24554=>X"00",
24555=>X"00",
24556=>X"00",
24557=>X"00",
24558=>X"00",
24559=>X"00",
24560=>X"00",
24561=>X"00",
24562=>X"00",
24563=>X"00",
24564=>X"00",
24565=>X"00",
24566=>X"00",
24567=>X"00",
24568=>X"00",
24569=>X"00",
24570=>X"00",
24571=>X"00",
24572=>X"00",
24573=>X"00",
24574=>X"00",
24575=>X"00",
24576=>X"00",
24577=>X"00",
24578=>X"00",
24579=>X"00",
24580=>X"00",
24581=>X"00",
24582=>X"00",
24583=>X"00",
24584=>X"00",
24585=>X"00",
24586=>X"00",
24587=>X"00",
24588=>X"00",
24589=>X"00",
24590=>X"00",
24591=>X"00",
24592=>X"00",
24593=>X"00",
24594=>X"00",
24595=>X"00",
24596=>X"00",
24597=>X"00",
24598=>X"00",
24599=>X"00",
24600=>X"00",
24601=>X"00",
24602=>X"00",
24603=>X"00",
24604=>X"00",
24605=>X"00",
24606=>X"00",
24607=>X"00",
24608=>X"00",
24609=>X"00",
24610=>X"00",
24611=>X"00",
24612=>X"00",
24613=>X"00",
24614=>X"00",
24615=>X"00",
24616=>X"00",
24617=>X"00",
24618=>X"00",
24619=>X"00",
24620=>X"00",
24621=>X"00",
24622=>X"00",
24623=>X"00",
24624=>X"00",
24625=>X"00",
24626=>X"00",
24627=>X"00",
24628=>X"00",
24629=>X"00",
24630=>X"00",
24631=>X"00",
24632=>X"00",
24633=>X"00",
24634=>X"00",
24635=>X"00",
24636=>X"00",
24637=>X"00",
24638=>X"00",
24639=>X"00",
24640=>X"00",
24641=>X"00",
24642=>X"00",
24643=>X"00",
24644=>X"00",
24645=>X"00",
24646=>X"00",
24647=>X"00",
24648=>X"00",
24649=>X"00",
24650=>X"00",
24651=>X"00",
24652=>X"00",
24653=>X"00",
24654=>X"00",
24655=>X"00",
24656=>X"00",
24657=>X"00",
24658=>X"00",
24659=>X"00",
24660=>X"00",
24661=>X"00",
24662=>X"00",
24663=>X"00",
24664=>X"00",
24665=>X"00",
24666=>X"00",
24667=>X"00",
24668=>X"00",
24669=>X"00",
24670=>X"00",
24671=>X"00",
24672=>X"00",
24673=>X"00",
24674=>X"00",
24675=>X"00",
24676=>X"00",
24677=>X"00",
24678=>X"00",
24679=>X"00",
24680=>X"00",
24681=>X"00",
24682=>X"00",
24683=>X"00",
24684=>X"00",
24685=>X"00",
24686=>X"00",
24687=>X"00",
24688=>X"00",
24689=>X"00",
24690=>X"00",
24691=>X"00",
24692=>X"00",
24693=>X"00",
24694=>X"00",
24695=>X"00",
24696=>X"00",
24697=>X"00",
24698=>X"00",
24699=>X"00",
24700=>X"00",
24701=>X"00",
24702=>X"00",
24703=>X"00",
24704=>X"00",
24705=>X"00",
24706=>X"00",
24707=>X"00",
24708=>X"00",
24709=>X"00",
24710=>X"00",
24711=>X"00",
24712=>X"00",
24713=>X"00",
24714=>X"00",
24715=>X"00",
24716=>X"00",
24717=>X"00",
24718=>X"00",
24719=>X"00",
24720=>X"00",
24721=>X"00",
24722=>X"00",
24723=>X"00",
24724=>X"00",
24725=>X"00",
24726=>X"00",
24727=>X"00",
24728=>X"00",
24729=>X"00",
24730=>X"00",
24731=>X"00",
24732=>X"00",
24733=>X"00",
24734=>X"00",
24735=>X"00",
24736=>X"00",
24737=>X"00",
24738=>X"00",
24739=>X"00",
24740=>X"00",
24741=>X"00",
24742=>X"00",
24743=>X"00",
24744=>X"00",
24745=>X"00",
24746=>X"00",
24747=>X"00",
24748=>X"00",
24749=>X"00",
24750=>X"00",
24751=>X"00",
24752=>X"00",
24753=>X"00",
24754=>X"00",
24755=>X"00",
24756=>X"00",
24757=>X"00",
24758=>X"00",
24759=>X"00",
24760=>X"00",
24761=>X"00",
24762=>X"00",
24763=>X"00",
24764=>X"00",
24765=>X"00",
24766=>X"00",
24767=>X"00",
24768=>X"00",
24769=>X"00",
24770=>X"00",
24771=>X"00",
24772=>X"00",
24773=>X"00",
24774=>X"00",
24775=>X"00",
24776=>X"00",
24777=>X"00",
24778=>X"00",
24779=>X"00",
24780=>X"00",
24781=>X"00",
24782=>X"00",
24783=>X"00",
24784=>X"00",
24785=>X"00",
24786=>X"00",
24787=>X"00",
24788=>X"00",
24789=>X"00",
24790=>X"00",
24791=>X"00",
24792=>X"00",
24793=>X"00",
24794=>X"00",
24795=>X"00",
24796=>X"00",
24797=>X"00",
24798=>X"00",
24799=>X"00",
24800=>X"00",
24801=>X"00",
24802=>X"00",
24803=>X"00",
24804=>X"00",
24805=>X"00",
24806=>X"00",
24807=>X"00",
24808=>X"00",
24809=>X"00",
24810=>X"00",
24811=>X"00",
24812=>X"00",
24813=>X"00",
24814=>X"00",
24815=>X"00",
24816=>X"00",
24817=>X"00",
24818=>X"00",
24819=>X"00",
24820=>X"00",
24821=>X"00",
24822=>X"00",
24823=>X"00",
24824=>X"00",
24825=>X"00",
24826=>X"00",
24827=>X"00",
24828=>X"00",
24829=>X"00",
24830=>X"00",
24831=>X"00",
24832=>X"00",
24833=>X"00",
24834=>X"00",
24835=>X"00",
24836=>X"00",
24837=>X"00",
24838=>X"00",
24839=>X"00",
24840=>X"00",
24841=>X"00",
24842=>X"00",
24843=>X"00",
24844=>X"00",
24845=>X"00",
24846=>X"00",
24847=>X"00",
24848=>X"00",
24849=>X"00",
24850=>X"00",
24851=>X"00",
24852=>X"00",
24853=>X"00",
24854=>X"00",
24855=>X"00",
24856=>X"00",
24857=>X"00",
24858=>X"00",
24859=>X"00",
24860=>X"00",
24861=>X"00",
24862=>X"00",
24863=>X"00",
24864=>X"00",
24865=>X"00",
24866=>X"00",
24867=>X"00",
24868=>X"00",
24869=>X"00",
24870=>X"00",
24871=>X"00",
24872=>X"00",
24873=>X"00",
24874=>X"00",
24875=>X"00",
24876=>X"00",
24877=>X"00",
24878=>X"00",
24879=>X"00",
24880=>X"00",
24881=>X"00",
24882=>X"00",
24883=>X"00",
24884=>X"00",
24885=>X"00",
24886=>X"00",
24887=>X"00",
24888=>X"00",
24889=>X"00",
24890=>X"00",
24891=>X"00",
24892=>X"00",
24893=>X"00",
24894=>X"00",
24895=>X"00",
24896=>X"00",
24897=>X"00",
24898=>X"00",
24899=>X"00",
24900=>X"00",
24901=>X"00",
24902=>X"00",
24903=>X"00",
24904=>X"00",
24905=>X"00",
24906=>X"00",
24907=>X"00",
24908=>X"00",
24909=>X"00",
24910=>X"00",
24911=>X"00",
24912=>X"00",
24913=>X"00",
24914=>X"00",
24915=>X"00",
24916=>X"00",
24917=>X"00",
24918=>X"00",
24919=>X"00",
24920=>X"00",
24921=>X"00",
24922=>X"00",
24923=>X"00",
24924=>X"00",
24925=>X"00",
24926=>X"00",
24927=>X"00",
24928=>X"00",
24929=>X"00",
24930=>X"00",
24931=>X"00",
24932=>X"00",
24933=>X"00",
24934=>X"00",
24935=>X"00",
24936=>X"00",
24937=>X"00",
24938=>X"00",
24939=>X"00",
24940=>X"00",
24941=>X"00",
24942=>X"00",
24943=>X"00",
24944=>X"00",
24945=>X"00",
24946=>X"00",
24947=>X"00",
24948=>X"00",
24949=>X"00",
24950=>X"00",
24951=>X"00",
24952=>X"00",
24953=>X"00",
24954=>X"00",
24955=>X"00",
24956=>X"00",
24957=>X"00",
24958=>X"00",
24959=>X"00",
24960=>X"00",
24961=>X"00",
24962=>X"00",
24963=>X"00",
24964=>X"00",
24965=>X"00",
24966=>X"00",
24967=>X"00",
24968=>X"00",
24969=>X"00",
24970=>X"00",
24971=>X"00",
24972=>X"00",
24973=>X"00",
24974=>X"00",
24975=>X"00",
24976=>X"00",
24977=>X"00",
24978=>X"00",
24979=>X"00",
24980=>X"00",
24981=>X"00",
24982=>X"00",
24983=>X"00",
24984=>X"00",
24985=>X"00",
24986=>X"00",
24987=>X"00",
24988=>X"00",
24989=>X"00",
24990=>X"00",
24991=>X"00",
24992=>X"00",
24993=>X"00",
24994=>X"00",
24995=>X"00",
24996=>X"00",
24997=>X"00",
24998=>X"00",
24999=>X"00",
25000=>X"00",
25001=>X"00",
25002=>X"00",
25003=>X"00",
25004=>X"00",
25005=>X"00",
25006=>X"00",
25007=>X"00",
25008=>X"00",
25009=>X"00",
25010=>X"00",
25011=>X"00",
25012=>X"00",
25013=>X"00",
25014=>X"00",
25015=>X"00",
25016=>X"00",
25017=>X"00",
25018=>X"00",
25019=>X"00",
25020=>X"00",
25021=>X"00",
25022=>X"00",
25023=>X"00",
25024=>X"00",
25025=>X"00",
25026=>X"00",
25027=>X"00",
25028=>X"00",
25029=>X"00",
25030=>X"00",
25031=>X"00",
25032=>X"00",
25033=>X"00",
25034=>X"00",
25035=>X"00",
25036=>X"00",
25037=>X"00",
25038=>X"00",
25039=>X"00",
25040=>X"00",
25041=>X"00",
25042=>X"00",
25043=>X"00",
25044=>X"00",
25045=>X"00",
25046=>X"00",
25047=>X"00",
25048=>X"00",
25049=>X"00",
25050=>X"00",
25051=>X"00",
25052=>X"00",
25053=>X"00",
25054=>X"00",
25055=>X"00",
25056=>X"00",
25057=>X"00",
25058=>X"00",
25059=>X"00",
25060=>X"00",
25061=>X"00",
25062=>X"00",
25063=>X"00",
25064=>X"00",
25065=>X"00",
25066=>X"00",
25067=>X"00",
25068=>X"00",
25069=>X"00",
25070=>X"00",
25071=>X"00",
25072=>X"00",
25073=>X"00",
25074=>X"00",
25075=>X"00",
25076=>X"00",
25077=>X"00",
25078=>X"00",
25079=>X"00",
25080=>X"00",
25081=>X"00",
25082=>X"00",
25083=>X"00",
25084=>X"00",
25085=>X"00",
25086=>X"00",
25087=>X"00",
25088=>X"00",
25089=>X"00",
25090=>X"00",
25091=>X"00",
25092=>X"00",
25093=>X"00",
25094=>X"00",
25095=>X"00",
25096=>X"00",
25097=>X"00",
25098=>X"00",
25099=>X"00",
25100=>X"00",
25101=>X"00",
25102=>X"00",
25103=>X"00",
25104=>X"00",
25105=>X"00",
25106=>X"00",
25107=>X"00",
25108=>X"00",
25109=>X"00",
25110=>X"00",
25111=>X"00",
25112=>X"00",
25113=>X"00",
25114=>X"00",
25115=>X"00",
25116=>X"00",
25117=>X"00",
25118=>X"00",
25119=>X"00",
25120=>X"00",
25121=>X"00",
25122=>X"00",
25123=>X"00",
25124=>X"00",
25125=>X"00",
25126=>X"00",
25127=>X"00",
25128=>X"00",
25129=>X"00",
25130=>X"00",
25131=>X"00",
25132=>X"00",
25133=>X"00",
25134=>X"00",
25135=>X"00",
25136=>X"00",
25137=>X"00",
25138=>X"00",
25139=>X"00",
25140=>X"00",
25141=>X"00",
25142=>X"00",
25143=>X"00",
25144=>X"00",
25145=>X"00",
25146=>X"00",
25147=>X"00",
25148=>X"00",
25149=>X"00",
25150=>X"00",
25151=>X"00",
25152=>X"00",
25153=>X"00",
25154=>X"00",
25155=>X"00",
25156=>X"00",
25157=>X"00",
25158=>X"00",
25159=>X"00",
25160=>X"00",
25161=>X"00",
25162=>X"00",
25163=>X"00",
25164=>X"00",
25165=>X"00",
25166=>X"00",
25167=>X"00",
25168=>X"00",
25169=>X"00",
25170=>X"00",
25171=>X"00",
25172=>X"00",
25173=>X"00",
25174=>X"00",
25175=>X"00",
25176=>X"00",
25177=>X"00",
25178=>X"00",
25179=>X"00",
25180=>X"00",
25181=>X"00",
25182=>X"00",
25183=>X"00",
25184=>X"00",
25185=>X"00",
25186=>X"00",
25187=>X"00",
25188=>X"00",
25189=>X"00",
25190=>X"00",
25191=>X"00",
25192=>X"00",
25193=>X"00",
25194=>X"00",
25195=>X"00",
25196=>X"00",
25197=>X"00",
25198=>X"00",
25199=>X"00",
25200=>X"00",
25201=>X"00",
25202=>X"00",
25203=>X"00",
25204=>X"00",
25205=>X"00",
25206=>X"00",
25207=>X"00",
25208=>X"00",
25209=>X"00",
25210=>X"00",
25211=>X"00",
25212=>X"00",
25213=>X"00",
25214=>X"00",
25215=>X"00",
25216=>X"00",
25217=>X"00",
25218=>X"00",
25219=>X"00",
25220=>X"00",
25221=>X"00",
25222=>X"00",
25223=>X"00",
25224=>X"00",
25225=>X"00",
25226=>X"00",
25227=>X"00",
25228=>X"00",
25229=>X"00",
25230=>X"00",
25231=>X"00",
25232=>X"00",
25233=>X"00",
25234=>X"00",
25235=>X"00",
25236=>X"00",
25237=>X"00",
25238=>X"00",
25239=>X"00",
25240=>X"00",
25241=>X"00",
25242=>X"00",
25243=>X"00",
25244=>X"00",
25245=>X"00",
25246=>X"00",
25247=>X"00",
25248=>X"00",
25249=>X"00",
25250=>X"00",
25251=>X"00",
25252=>X"00",
25253=>X"00",
25254=>X"00",
25255=>X"00",
25256=>X"00",
25257=>X"00",
25258=>X"00",
25259=>X"00",
25260=>X"00",
25261=>X"00",
25262=>X"00",
25263=>X"00",
25264=>X"00",
25265=>X"00",
25266=>X"00",
25267=>X"00",
25268=>X"00",
25269=>X"00",
25270=>X"00",
25271=>X"00",
25272=>X"00",
25273=>X"00",
25274=>X"00",
25275=>X"00",
25276=>X"00",
25277=>X"00",
25278=>X"00",
25279=>X"00",
25280=>X"00",
25281=>X"00",
25282=>X"00",
25283=>X"00",
25284=>X"00",
25285=>X"00",
25286=>X"00",
25287=>X"00",
25288=>X"00",
25289=>X"00",
25290=>X"00",
25291=>X"00",
25292=>X"00",
25293=>X"00",
25294=>X"00",
25295=>X"00",
25296=>X"00",
25297=>X"00",
25298=>X"00",
25299=>X"00",
25300=>X"00",
25301=>X"00",
25302=>X"00",
25303=>X"00",
25304=>X"00",
25305=>X"00",
25306=>X"00",
25307=>X"00",
25308=>X"00",
25309=>X"00",
25310=>X"00",
25311=>X"00",
25312=>X"00",
25313=>X"00",
25314=>X"00",
25315=>X"00",
25316=>X"00",
25317=>X"00",
25318=>X"00",
25319=>X"00",
25320=>X"00",
25321=>X"00",
25322=>X"00",
25323=>X"00",
25324=>X"00",
25325=>X"00",
25326=>X"00",
25327=>X"00",
25328=>X"00",
25329=>X"00",
25330=>X"00",
25331=>X"00",
25332=>X"00",
25333=>X"00",
25334=>X"00",
25335=>X"00",
25336=>X"00",
25337=>X"00",
25338=>X"00",
25339=>X"00",
25340=>X"00",
25341=>X"00",
25342=>X"00",
25343=>X"00",
25344=>X"00",
25345=>X"00",
25346=>X"00",
25347=>X"00",
25348=>X"00",
25349=>X"00",
25350=>X"00",
25351=>X"00",
25352=>X"00",
25353=>X"00",
25354=>X"00",
25355=>X"00",
25356=>X"00",
25357=>X"00",
25358=>X"00",
25359=>X"00",
25360=>X"00",
25361=>X"00",
25362=>X"00",
25363=>X"00",
25364=>X"00",
25365=>X"00",
25366=>X"00",
25367=>X"00",
25368=>X"00",
25369=>X"00",
25370=>X"00",
25371=>X"00",
25372=>X"00",
25373=>X"00",
25374=>X"00",
25375=>X"00",
25376=>X"00",
25377=>X"00",
25378=>X"00",
25379=>X"00",
25380=>X"00",
25381=>X"00",
25382=>X"00",
25383=>X"00",
25384=>X"00",
25385=>X"00",
25386=>X"00",
25387=>X"00",
25388=>X"00",
25389=>X"00",
25390=>X"00",
25391=>X"00",
25392=>X"00",
25393=>X"00",
25394=>X"00",
25395=>X"00",
25396=>X"00",
25397=>X"00",
25398=>X"00",
25399=>X"00",
25400=>X"00",
25401=>X"00",
25402=>X"00",
25403=>X"00",
25404=>X"00",
25405=>X"00",
25406=>X"00",
25407=>X"00",
25408=>X"00",
25409=>X"00",
25410=>X"00",
25411=>X"00",
25412=>X"00",
25413=>X"00",
25414=>X"00",
25415=>X"00",
25416=>X"00",
25417=>X"00",
25418=>X"00",
25419=>X"00",
25420=>X"00",
25421=>X"00",
25422=>X"00",
25423=>X"00",
25424=>X"00",
25425=>X"00",
25426=>X"00",
25427=>X"00",
25428=>X"00",
25429=>X"00",
25430=>X"00",
25431=>X"00",
25432=>X"00",
25433=>X"00",
25434=>X"00",
25435=>X"00",
25436=>X"00",
25437=>X"00",
25438=>X"00",
25439=>X"00",
25440=>X"00",
25441=>X"00",
25442=>X"00",
25443=>X"00",
25444=>X"00",
25445=>X"00",
25446=>X"00",
25447=>X"00",
25448=>X"00",
25449=>X"00",
25450=>X"00",
25451=>X"00",
25452=>X"00",
25453=>X"00",
25454=>X"00",
25455=>X"00",
25456=>X"00",
25457=>X"00",
25458=>X"00",
25459=>X"00",
25460=>X"00",
25461=>X"00",
25462=>X"00",
25463=>X"00",
25464=>X"00",
25465=>X"00",
25466=>X"00",
25467=>X"00",
25468=>X"00",
25469=>X"00",
25470=>X"00",
25471=>X"00",
25472=>X"00",
25473=>X"00",
25474=>X"00",
25475=>X"00",
25476=>X"00",
25477=>X"00",
25478=>X"00",
25479=>X"00",
25480=>X"00",
25481=>X"00",
25482=>X"00",
25483=>X"00",
25484=>X"00",
25485=>X"00",
25486=>X"00",
25487=>X"00",
25488=>X"00",
25489=>X"00",
25490=>X"00",
25491=>X"00",
25492=>X"00",
25493=>X"00",
25494=>X"00",
25495=>X"00",
25496=>X"00",
25497=>X"00",
25498=>X"00",
25499=>X"00",
25500=>X"00",
25501=>X"00",
25502=>X"00",
25503=>X"00",
25504=>X"00",
25505=>X"00",
25506=>X"00",
25507=>X"00",
25508=>X"00",
25509=>X"00",
25510=>X"00",
25511=>X"00",
25512=>X"00",
25513=>X"00",
25514=>X"00",
25515=>X"00",
25516=>X"00",
25517=>X"00",
25518=>X"00",
25519=>X"00",
25520=>X"00",
25521=>X"00",
25522=>X"00",
25523=>X"00",
25524=>X"00",
25525=>X"00",
25526=>X"00",
25527=>X"00",
25528=>X"00",
25529=>X"00",
25530=>X"00",
25531=>X"00",
25532=>X"00",
25533=>X"00",
25534=>X"00",
25535=>X"00",
25536=>X"00",
25537=>X"00",
25538=>X"00",
25539=>X"00",
25540=>X"00",
25541=>X"00",
25542=>X"00",
25543=>X"00",
25544=>X"00",
25545=>X"00",
25546=>X"00",
25547=>X"00",
25548=>X"00",
25549=>X"00",
25550=>X"00",
25551=>X"00",
25552=>X"00",
25553=>X"00",
25554=>X"00",
25555=>X"00",
25556=>X"00",
25557=>X"00",
25558=>X"00",
25559=>X"00",
25560=>X"00",
25561=>X"00",
25562=>X"00",
25563=>X"00",
25564=>X"00",
25565=>X"00",
25566=>X"00",
25567=>X"00",
25568=>X"00",
25569=>X"00",
25570=>X"00",
25571=>X"00",
25572=>X"00",
25573=>X"00",
25574=>X"00",
25575=>X"00",
25576=>X"00",
25577=>X"00",
25578=>X"00",
25579=>X"00",
25580=>X"00",
25581=>X"00",
25582=>X"00",
25583=>X"00",
25584=>X"00",
25585=>X"00",
25586=>X"00",
25587=>X"00",
25588=>X"00",
25589=>X"00",
25590=>X"00",
25591=>X"00",
25592=>X"00",
25593=>X"00",
25594=>X"00",
25595=>X"00",
25596=>X"00",
25597=>X"00",
25598=>X"00",
25599=>X"00",
25600=>X"00",
25601=>X"00",
25602=>X"00",
25603=>X"00",
25604=>X"00",
25605=>X"00",
25606=>X"00",
25607=>X"00",
25608=>X"00",
25609=>X"00",
25610=>X"00",
25611=>X"00",
25612=>X"00",
25613=>X"00",
25614=>X"00",
25615=>X"00",
25616=>X"00",
25617=>X"00",
25618=>X"00",
25619=>X"00",
25620=>X"00",
25621=>X"00",
25622=>X"00",
25623=>X"00",
25624=>X"00",
25625=>X"00",
25626=>X"00",
25627=>X"00",
25628=>X"00",
25629=>X"00",
25630=>X"00",
25631=>X"00",
25632=>X"00",
25633=>X"00",
25634=>X"00",
25635=>X"00",
25636=>X"00",
25637=>X"00",
25638=>X"00",
25639=>X"00",
25640=>X"00",
25641=>X"00",
25642=>X"00",
25643=>X"00",
25644=>X"00",
25645=>X"00",
25646=>X"00",
25647=>X"00",
25648=>X"00",
25649=>X"00",
25650=>X"00",
25651=>X"00",
25652=>X"00",
25653=>X"00",
25654=>X"00",
25655=>X"00",
25656=>X"00",
25657=>X"00",
25658=>X"00",
25659=>X"00",
25660=>X"00",
25661=>X"00",
25662=>X"00",
25663=>X"00",
25664=>X"00",
25665=>X"00",
25666=>X"00",
25667=>X"00",
25668=>X"00",
25669=>X"00",
25670=>X"00",
25671=>X"00",
25672=>X"00",
25673=>X"00",
25674=>X"00",
25675=>X"00",
25676=>X"00",
25677=>X"00",
25678=>X"00",
25679=>X"00",
25680=>X"00",
25681=>X"00",
25682=>X"00",
25683=>X"00",
25684=>X"00",
25685=>X"00",
25686=>X"00",
25687=>X"00",
25688=>X"00",
25689=>X"00",
25690=>X"00",
25691=>X"00",
25692=>X"00",
25693=>X"00",
25694=>X"00",
25695=>X"00",
25696=>X"00",
25697=>X"00",
25698=>X"00",
25699=>X"00",
25700=>X"00",
25701=>X"00",
25702=>X"00",
25703=>X"00",
25704=>X"00",
25705=>X"00",
25706=>X"00",
25707=>X"00",
25708=>X"00",
25709=>X"00",
25710=>X"00",
25711=>X"00",
25712=>X"00",
25713=>X"00",
25714=>X"00",
25715=>X"00",
25716=>X"00",
25717=>X"00",
25718=>X"00",
25719=>X"00",
25720=>X"00",
25721=>X"00",
25722=>X"00",
25723=>X"00",
25724=>X"00",
25725=>X"00",
25726=>X"00",
25727=>X"00",
25728=>X"00",
25729=>X"00",
25730=>X"00",
25731=>X"00",
25732=>X"00",
25733=>X"00",
25734=>X"00",
25735=>X"00",
25736=>X"00",
25737=>X"00",
25738=>X"00",
25739=>X"00",
25740=>X"00",
25741=>X"00",
25742=>X"00",
25743=>X"00",
25744=>X"00",
25745=>X"00",
25746=>X"00",
25747=>X"00",
25748=>X"00",
25749=>X"00",
25750=>X"00",
25751=>X"00",
25752=>X"00",
25753=>X"00",
25754=>X"00",
25755=>X"00",
25756=>X"00",
25757=>X"00",
25758=>X"00",
25759=>X"00",
25760=>X"00",
25761=>X"00",
25762=>X"00",
25763=>X"00",
25764=>X"00",
25765=>X"00",
25766=>X"00",
25767=>X"00",
25768=>X"00",
25769=>X"00",
25770=>X"00",
25771=>X"00",
25772=>X"00",
25773=>X"00",
25774=>X"00",
25775=>X"00",
25776=>X"00",
25777=>X"00",
25778=>X"00",
25779=>X"00",
25780=>X"00",
25781=>X"00",
25782=>X"00",
25783=>X"00",
25784=>X"00",
25785=>X"00",
25786=>X"00",
25787=>X"00",
25788=>X"00",
25789=>X"00",
25790=>X"00",
25791=>X"00",
25792=>X"00",
25793=>X"00",
25794=>X"00",
25795=>X"00",
25796=>X"00",
25797=>X"00",
25798=>X"00",
25799=>X"00",
25800=>X"00",
25801=>X"00",
25802=>X"00",
25803=>X"00",
25804=>X"00",
25805=>X"00",
25806=>X"00",
25807=>X"00",
25808=>X"00",
25809=>X"00",
25810=>X"00",
25811=>X"00",
25812=>X"00",
25813=>X"00",
25814=>X"00",
25815=>X"00",
25816=>X"00",
25817=>X"00",
25818=>X"00",
25819=>X"00",
25820=>X"00",
25821=>X"00",
25822=>X"00",
25823=>X"00",
25824=>X"00",
25825=>X"00",
25826=>X"00",
25827=>X"00",
25828=>X"00",
25829=>X"00",
25830=>X"00",
25831=>X"00",
25832=>X"00",
25833=>X"00",
25834=>X"00",
25835=>X"00",
25836=>X"00",
25837=>X"00",
25838=>X"00",
25839=>X"00",
25840=>X"00",
25841=>X"00",
25842=>X"00",
25843=>X"00",
25844=>X"00",
25845=>X"00",
25846=>X"00",
25847=>X"00",
25848=>X"00",
25849=>X"00",
25850=>X"00",
25851=>X"00",
25852=>X"00",
25853=>X"00",
25854=>X"00",
25855=>X"00",
25856=>X"00",
25857=>X"00",
25858=>X"00",
25859=>X"00",
25860=>X"00",
25861=>X"00",
25862=>X"00",
25863=>X"00",
25864=>X"00",
25865=>X"00",
25866=>X"00",
25867=>X"00",
25868=>X"00",
25869=>X"00",
25870=>X"00",
25871=>X"00",
25872=>X"00",
25873=>X"00",
25874=>X"00",
25875=>X"00",
25876=>X"00",
25877=>X"00",
25878=>X"00",
25879=>X"00",
25880=>X"00",
25881=>X"00",
25882=>X"00",
25883=>X"00",
25884=>X"00",
25885=>X"00",
25886=>X"00",
25887=>X"00",
25888=>X"00",
25889=>X"00",
25890=>X"00",
25891=>X"00",
25892=>X"00",
25893=>X"00",
25894=>X"00",
25895=>X"00",
25896=>X"00",
25897=>X"00",
25898=>X"00",
25899=>X"00",
25900=>X"00",
25901=>X"00",
25902=>X"00",
25903=>X"00",
25904=>X"00",
25905=>X"00",
25906=>X"00",
25907=>X"00",
25908=>X"00",
25909=>X"00",
25910=>X"00",
25911=>X"00",
25912=>X"00",
25913=>X"00",
25914=>X"00",
25915=>X"00",
25916=>X"00",
25917=>X"00",
25918=>X"00",
25919=>X"00",
25920=>X"00",
25921=>X"00",
25922=>X"00",
25923=>X"00",
25924=>X"00",
25925=>X"00",
25926=>X"00",
25927=>X"00",
25928=>X"00",
25929=>X"00",
25930=>X"00",
25931=>X"00",
25932=>X"00",
25933=>X"00",
25934=>X"00",
25935=>X"00",
25936=>X"00",
25937=>X"00",
25938=>X"00",
25939=>X"00",
25940=>X"00",
25941=>X"00",
25942=>X"00",
25943=>X"00",
25944=>X"00",
25945=>X"00",
25946=>X"00",
25947=>X"00",
25948=>X"00",
25949=>X"00",
25950=>X"00",
25951=>X"00",
25952=>X"00",
25953=>X"00",
25954=>X"00",
25955=>X"00",
25956=>X"00",
25957=>X"00",
25958=>X"00",
25959=>X"00",
25960=>X"00",
25961=>X"00",
25962=>X"00",
25963=>X"00",
25964=>X"00",
25965=>X"00",
25966=>X"00",
25967=>X"00",
25968=>X"00",
25969=>X"00",
25970=>X"00",
25971=>X"00",
25972=>X"00",
25973=>X"00",
25974=>X"00",
25975=>X"00",
25976=>X"00",
25977=>X"00",
25978=>X"00",
25979=>X"00",
25980=>X"00",
25981=>X"00",
25982=>X"00",
25983=>X"00",
25984=>X"00",
25985=>X"00",
25986=>X"00",
25987=>X"00",
25988=>X"00",
25989=>X"00",
25990=>X"00",
25991=>X"00",
25992=>X"00",
25993=>X"00",
25994=>X"00",
25995=>X"00",
25996=>X"00",
25997=>X"00",
25998=>X"00",
25999=>X"00",
26000=>X"00",
26001=>X"00",
26002=>X"00",
26003=>X"00",
26004=>X"00",
26005=>X"00",
26006=>X"00",
26007=>X"00",
26008=>X"00",
26009=>X"00",
26010=>X"00",
26011=>X"00",
26012=>X"00",
26013=>X"00",
26014=>X"00",
26015=>X"00",
26016=>X"00",
26017=>X"00",
26018=>X"00",
26019=>X"00",
26020=>X"00",
26021=>X"00",
26022=>X"00",
26023=>X"00",
26024=>X"00",
26025=>X"00",
26026=>X"00",
26027=>X"00",
26028=>X"00",
26029=>X"00",
26030=>X"00",
26031=>X"00",
26032=>X"00",
26033=>X"00",
26034=>X"00",
26035=>X"00",
26036=>X"00",
26037=>X"00",
26038=>X"00",
26039=>X"00",
26040=>X"00",
26041=>X"00",
26042=>X"00",
26043=>X"00",
26044=>X"00",
26045=>X"00",
26046=>X"00",
26047=>X"00",
26048=>X"00",
26049=>X"00",
26050=>X"00",
26051=>X"00",
26052=>X"00",
26053=>X"00",
26054=>X"00",
26055=>X"00",
26056=>X"00",
26057=>X"00",
26058=>X"00",
26059=>X"00",
26060=>X"00",
26061=>X"00",
26062=>X"00",
26063=>X"00",
26064=>X"00",
26065=>X"00",
26066=>X"00",
26067=>X"00",
26068=>X"00",
26069=>X"00",
26070=>X"00",
26071=>X"00",
26072=>X"00",
26073=>X"00",
26074=>X"00",
26075=>X"00",
26076=>X"00",
26077=>X"00",
26078=>X"00",
26079=>X"00",
26080=>X"00",
26081=>X"00",
26082=>X"00",
26083=>X"00",
26084=>X"00",
26085=>X"00",
26086=>X"00",
26087=>X"00",
26088=>X"00",
26089=>X"00",
26090=>X"00",
26091=>X"00",
26092=>X"00",
26093=>X"00",
26094=>X"00",
26095=>X"00",
26096=>X"00",
26097=>X"00",
26098=>X"00",
26099=>X"00",
26100=>X"00",
26101=>X"00",
26102=>X"00",
26103=>X"00",
26104=>X"00",
26105=>X"00",
26106=>X"00",
26107=>X"00",
26108=>X"00",
26109=>X"00",
26110=>X"00",
26111=>X"00",
26112=>X"00",
26113=>X"00",
26114=>X"00",
26115=>X"00",
26116=>X"00",
26117=>X"00",
26118=>X"00",
26119=>X"00",
26120=>X"00",
26121=>X"00",
26122=>X"00",
26123=>X"00",
26124=>X"00",
26125=>X"00",
26126=>X"00",
26127=>X"00",
26128=>X"00",
26129=>X"00",
26130=>X"00",
26131=>X"00",
26132=>X"00",
26133=>X"00",
26134=>X"00",
26135=>X"00",
26136=>X"00",
26137=>X"00",
26138=>X"00",
26139=>X"00",
26140=>X"00",
26141=>X"00",
26142=>X"00",
26143=>X"00",
26144=>X"00",
26145=>X"00",
26146=>X"00",
26147=>X"00",
26148=>X"00",
26149=>X"00",
26150=>X"00",
26151=>X"00",
26152=>X"00",
26153=>X"00",
26154=>X"00",
26155=>X"00",
26156=>X"00",
26157=>X"00",
26158=>X"00",
26159=>X"00",
26160=>X"00",
26161=>X"00",
26162=>X"00",
26163=>X"00",
26164=>X"00",
26165=>X"00",
26166=>X"00",
26167=>X"00",
26168=>X"00",
26169=>X"00",
26170=>X"00",
26171=>X"00",
26172=>X"00",
26173=>X"00",
26174=>X"00",
26175=>X"00",
26176=>X"00",
26177=>X"00",
26178=>X"00",
26179=>X"00",
26180=>X"00",
26181=>X"00",
26182=>X"00",
26183=>X"00",
26184=>X"00",
26185=>X"00",
26186=>X"00",
26187=>X"00",
26188=>X"00",
26189=>X"00",
26190=>X"00",
26191=>X"00",
26192=>X"00",
26193=>X"00",
26194=>X"00",
26195=>X"00",
26196=>X"00",
26197=>X"00",
26198=>X"00",
26199=>X"00",
26200=>X"00",
26201=>X"00",
26202=>X"00",
26203=>X"00",
26204=>X"00",
26205=>X"00",
26206=>X"00",
26207=>X"00",
26208=>X"00",
26209=>X"00",
26210=>X"00",
26211=>X"00",
26212=>X"00",
26213=>X"00",
26214=>X"00",
26215=>X"00",
26216=>X"00",
26217=>X"00",
26218=>X"00",
26219=>X"00",
26220=>X"00",
26221=>X"00",
26222=>X"00",
26223=>X"00",
26224=>X"00",
26225=>X"00",
26226=>X"00",
26227=>X"00",
26228=>X"00",
26229=>X"00",
26230=>X"00",
26231=>X"00",
26232=>X"00",
26233=>X"00",
26234=>X"00",
26235=>X"00",
26236=>X"00",
26237=>X"00",
26238=>X"00",
26239=>X"00",
26240=>X"00",
26241=>X"00",
26242=>X"00",
26243=>X"00",
26244=>X"00",
26245=>X"00",
26246=>X"00",
26247=>X"00",
26248=>X"00",
26249=>X"00",
26250=>X"00",
26251=>X"00",
26252=>X"00",
26253=>X"00",
26254=>X"00",
26255=>X"00",
26256=>X"00",
26257=>X"00",
26258=>X"00",
26259=>X"00",
26260=>X"00",
26261=>X"00",
26262=>X"00",
26263=>X"00",
26264=>X"00",
26265=>X"00",
26266=>X"00",
26267=>X"00",
26268=>X"00",
26269=>X"00",
26270=>X"00",
26271=>X"00",
26272=>X"00",
26273=>X"00",
26274=>X"00",
26275=>X"00",
26276=>X"00",
26277=>X"00",
26278=>X"00",
26279=>X"00",
26280=>X"00",
26281=>X"00",
26282=>X"00",
26283=>X"00",
26284=>X"00",
26285=>X"00",
26286=>X"00",
26287=>X"00",
26288=>X"00",
26289=>X"00",
26290=>X"00",
26291=>X"00",
26292=>X"00",
26293=>X"00",
26294=>X"00",
26295=>X"00",
26296=>X"00",
26297=>X"00",
26298=>X"00",
26299=>X"00",
26300=>X"00",
26301=>X"00",
26302=>X"00",
26303=>X"00",
26304=>X"00",
26305=>X"00",
26306=>X"00",
26307=>X"00",
26308=>X"00",
26309=>X"00",
26310=>X"00",
26311=>X"00",
26312=>X"00",
26313=>X"00",
26314=>X"00",
26315=>X"00",
26316=>X"00",
26317=>X"00",
26318=>X"00",
26319=>X"00",
26320=>X"00",
26321=>X"00",
26322=>X"00",
26323=>X"00",
26324=>X"00",
26325=>X"00",
26326=>X"00",
26327=>X"00",
26328=>X"00",
26329=>X"00",
26330=>X"00",
26331=>X"00",
26332=>X"00",
26333=>X"00",
26334=>X"00",
26335=>X"00",
26336=>X"00",
26337=>X"00",
26338=>X"00",
26339=>X"00",
26340=>X"00",
26341=>X"00",
26342=>X"00",
26343=>X"00",
26344=>X"00",
26345=>X"00",
26346=>X"00",
26347=>X"00",
26348=>X"00",
26349=>X"00",
26350=>X"00",
26351=>X"00",
26352=>X"00",
26353=>X"00",
26354=>X"00",
26355=>X"00",
26356=>X"00",
26357=>X"00",
26358=>X"00",
26359=>X"00",
26360=>X"00",
26361=>X"00",
26362=>X"00",
26363=>X"00",
26364=>X"00",
26365=>X"00",
26366=>X"00",
26367=>X"00",
26368=>X"00",
26369=>X"00",
26370=>X"00",
26371=>X"00",
26372=>X"00",
26373=>X"00",
26374=>X"00",
26375=>X"00",
26376=>X"00",
26377=>X"00",
26378=>X"00",
26379=>X"00",
26380=>X"00",
26381=>X"00",
26382=>X"00",
26383=>X"00",
26384=>X"00",
26385=>X"00",
26386=>X"00",
26387=>X"00",
26388=>X"00",
26389=>X"00",
26390=>X"00",
26391=>X"00",
26392=>X"00",
26393=>X"00",
26394=>X"00",
26395=>X"00",
26396=>X"00",
26397=>X"00",
26398=>X"00",
26399=>X"00",
26400=>X"00",
26401=>X"00",
26402=>X"00",
26403=>X"00",
26404=>X"00",
26405=>X"00",
26406=>X"00",
26407=>X"00",
26408=>X"00",
26409=>X"00",
26410=>X"00",
26411=>X"00",
26412=>X"00",
26413=>X"00",
26414=>X"00",
26415=>X"00",
26416=>X"00",
26417=>X"00",
26418=>X"00",
26419=>X"00",
26420=>X"00",
26421=>X"00",
26422=>X"00",
26423=>X"00",
26424=>X"00",
26425=>X"00",
26426=>X"00",
26427=>X"00",
26428=>X"00",
26429=>X"00",
26430=>X"00",
26431=>X"00",
26432=>X"00",
26433=>X"00",
26434=>X"00",
26435=>X"00",
26436=>X"00",
26437=>X"00",
26438=>X"00",
26439=>X"00",
26440=>X"00",
26441=>X"00",
26442=>X"00",
26443=>X"00",
26444=>X"00",
26445=>X"00",
26446=>X"00",
26447=>X"00",
26448=>X"00",
26449=>X"00",
26450=>X"00",
26451=>X"00",
26452=>X"00",
26453=>X"00",
26454=>X"00",
26455=>X"00",
26456=>X"00",
26457=>X"00",
26458=>X"00",
26459=>X"00",
26460=>X"00",
26461=>X"00",
26462=>X"00",
26463=>X"00",
26464=>X"00",
26465=>X"00",
26466=>X"00",
26467=>X"00",
26468=>X"00",
26469=>X"00",
26470=>X"00",
26471=>X"00",
26472=>X"00",
26473=>X"00",
26474=>X"00",
26475=>X"00",
26476=>X"00",
26477=>X"00",
26478=>X"00",
26479=>X"00",
26480=>X"00",
26481=>X"00",
26482=>X"00",
26483=>X"00",
26484=>X"00",
26485=>X"00",
26486=>X"00",
26487=>X"00",
26488=>X"00",
26489=>X"00",
26490=>X"00",
26491=>X"00",
26492=>X"00",
26493=>X"00",
26494=>X"00",
26495=>X"00",
26496=>X"00",
26497=>X"00",
26498=>X"00",
26499=>X"00",
26500=>X"00",
26501=>X"00",
26502=>X"00",
26503=>X"00",
26504=>X"00",
26505=>X"00",
26506=>X"00",
26507=>X"00",
26508=>X"00",
26509=>X"00",
26510=>X"00",
26511=>X"00",
26512=>X"00",
26513=>X"00",
26514=>X"00",
26515=>X"00",
26516=>X"00",
26517=>X"00",
26518=>X"00",
26519=>X"00",
26520=>X"00",
26521=>X"00",
26522=>X"00",
26523=>X"00",
26524=>X"00",
26525=>X"00",
26526=>X"00",
26527=>X"00",
26528=>X"00",
26529=>X"00",
26530=>X"00",
26531=>X"00",
26532=>X"00",
26533=>X"00",
26534=>X"00",
26535=>X"00",
26536=>X"00",
26537=>X"00",
26538=>X"00",
26539=>X"00",
26540=>X"00",
26541=>X"00",
26542=>X"00",
26543=>X"00",
26544=>X"00",
26545=>X"00",
26546=>X"00",
26547=>X"00",
26548=>X"00",
26549=>X"00",
26550=>X"00",
26551=>X"00",
26552=>X"00",
26553=>X"00",
26554=>X"00",
26555=>X"00",
26556=>X"00",
26557=>X"00",
26558=>X"00",
26559=>X"00",
26560=>X"00",
26561=>X"00",
26562=>X"00",
26563=>X"00",
26564=>X"00",
26565=>X"00",
26566=>X"00",
26567=>X"00",
26568=>X"00",
26569=>X"00",
26570=>X"00",
26571=>X"00",
26572=>X"00",
26573=>X"00",
26574=>X"00",
26575=>X"00",
26576=>X"00",
26577=>X"00",
26578=>X"00",
26579=>X"00",
26580=>X"00",
26581=>X"00",
26582=>X"00",
26583=>X"00",
26584=>X"00",
26585=>X"00",
26586=>X"00",
26587=>X"00",
26588=>X"00",
26589=>X"00",
26590=>X"00",
26591=>X"00",
26592=>X"00",
26593=>X"00",
26594=>X"00",
26595=>X"00",
26596=>X"00",
26597=>X"00",
26598=>X"00",
26599=>X"00",
26600=>X"00",
26601=>X"00",
26602=>X"00",
26603=>X"00",
26604=>X"00",
26605=>X"00",
26606=>X"00",
26607=>X"00",
26608=>X"00",
26609=>X"00",
26610=>X"00",
26611=>X"00",
26612=>X"00",
26613=>X"00",
26614=>X"00",
26615=>X"00",
26616=>X"00",
26617=>X"00",
26618=>X"00",
26619=>X"00",
26620=>X"00",
26621=>X"00",
26622=>X"00",
26623=>X"00",
26624=>X"00",
26625=>X"00",
26626=>X"00",
26627=>X"00",
26628=>X"00",
26629=>X"00",
26630=>X"00",
26631=>X"00",
26632=>X"00",
26633=>X"00",
26634=>X"00",
26635=>X"00",
26636=>X"00",
26637=>X"00",
26638=>X"00",
26639=>X"00",
26640=>X"00",
26641=>X"00",
26642=>X"00",
26643=>X"00",
26644=>X"00",
26645=>X"00",
26646=>X"00",
26647=>X"00",
26648=>X"00",
26649=>X"00",
26650=>X"00",
26651=>X"00",
26652=>X"00",
26653=>X"00",
26654=>X"00",
26655=>X"00",
26656=>X"00",
26657=>X"00",
26658=>X"00",
26659=>X"00",
26660=>X"00",
26661=>X"00",
26662=>X"00",
26663=>X"00",
26664=>X"00",
26665=>X"00",
26666=>X"00",
26667=>X"00",
26668=>X"00",
26669=>X"00",
26670=>X"00",
26671=>X"00",
26672=>X"00",
26673=>X"00",
26674=>X"00",
26675=>X"00",
26676=>X"00",
26677=>X"00",
26678=>X"00",
26679=>X"00",
26680=>X"00",
26681=>X"00",
26682=>X"00",
26683=>X"00",
26684=>X"00",
26685=>X"00",
26686=>X"00",
26687=>X"00",
26688=>X"00",
26689=>X"00",
26690=>X"00",
26691=>X"00",
26692=>X"00",
26693=>X"00",
26694=>X"00",
26695=>X"00",
26696=>X"00",
26697=>X"00",
26698=>X"00",
26699=>X"00",
26700=>X"00",
26701=>X"00",
26702=>X"00",
26703=>X"00",
26704=>X"00",
26705=>X"00",
26706=>X"00",
26707=>X"00",
26708=>X"00",
26709=>X"00",
26710=>X"00",
26711=>X"00",
26712=>X"00",
26713=>X"00",
26714=>X"00",
26715=>X"00",
26716=>X"00",
26717=>X"00",
26718=>X"00",
26719=>X"00",
26720=>X"00",
26721=>X"00",
26722=>X"00",
26723=>X"00",
26724=>X"00",
26725=>X"00",
26726=>X"00",
26727=>X"00",
26728=>X"00",
26729=>X"00",
26730=>X"00",
26731=>X"00",
26732=>X"00",
26733=>X"00",
26734=>X"00",
26735=>X"00",
26736=>X"00",
26737=>X"00",
26738=>X"00",
26739=>X"00",
26740=>X"00",
26741=>X"00",
26742=>X"00",
26743=>X"00",
26744=>X"00",
26745=>X"00",
26746=>X"00",
26747=>X"00",
26748=>X"00",
26749=>X"00",
26750=>X"00",
26751=>X"00",
26752=>X"00",
26753=>X"00",
26754=>X"00",
26755=>X"00",
26756=>X"00",
26757=>X"00",
26758=>X"00",
26759=>X"00",
26760=>X"00",
26761=>X"00",
26762=>X"00",
26763=>X"00",
26764=>X"00",
26765=>X"00",
26766=>X"00",
26767=>X"00",
26768=>X"00",
26769=>X"00",
26770=>X"00",
26771=>X"00",
26772=>X"00",
26773=>X"00",
26774=>X"00",
26775=>X"00",
26776=>X"00",
26777=>X"00",
26778=>X"00",
26779=>X"00",
26780=>X"00",
26781=>X"00",
26782=>X"00",
26783=>X"00",
26784=>X"00",
26785=>X"00",
26786=>X"00",
26787=>X"00",
26788=>X"00",
26789=>X"00",
26790=>X"00",
26791=>X"00",
26792=>X"00",
26793=>X"00",
26794=>X"00",
26795=>X"00",
26796=>X"00",
26797=>X"00",
26798=>X"00",
26799=>X"00",
26800=>X"00",
26801=>X"00",
26802=>X"00",
26803=>X"00",
26804=>X"00",
26805=>X"00",
26806=>X"00",
26807=>X"00",
26808=>X"00",
26809=>X"00",
26810=>X"00",
26811=>X"00",
26812=>X"00",
26813=>X"00",
26814=>X"00",
26815=>X"00",
26816=>X"00",
26817=>X"00",
26818=>X"00",
26819=>X"00",
26820=>X"00",
26821=>X"00",
26822=>X"00",
26823=>X"00",
26824=>X"00",
26825=>X"00",
26826=>X"00",
26827=>X"00",
26828=>X"00",
26829=>X"00",
26830=>X"00",
26831=>X"00",
26832=>X"00",
26833=>X"00",
26834=>X"00",
26835=>X"00",
26836=>X"00",
26837=>X"00",
26838=>X"00",
26839=>X"00",
26840=>X"00",
26841=>X"00",
26842=>X"00",
26843=>X"00",
26844=>X"00",
26845=>X"00",
26846=>X"00",
26847=>X"00",
26848=>X"00",
26849=>X"00",
26850=>X"00",
26851=>X"00",
26852=>X"00",
26853=>X"00",
26854=>X"00",
26855=>X"00",
26856=>X"00",
26857=>X"00",
26858=>X"00",
26859=>X"00",
26860=>X"00",
26861=>X"00",
26862=>X"00",
26863=>X"00",
26864=>X"00",
26865=>X"00",
26866=>X"00",
26867=>X"00",
26868=>X"00",
26869=>X"00",
26870=>X"00",
26871=>X"00",
26872=>X"00",
26873=>X"00",
26874=>X"00",
26875=>X"00",
26876=>X"00",
26877=>X"00",
26878=>X"00",
26879=>X"00",
26880=>X"00",
26881=>X"00",
26882=>X"00",
26883=>X"00",
26884=>X"00",
26885=>X"00",
26886=>X"00",
26887=>X"00",
26888=>X"00",
26889=>X"00",
26890=>X"00",
26891=>X"00",
26892=>X"00",
26893=>X"00",
26894=>X"00",
26895=>X"00",
26896=>X"00",
26897=>X"00",
26898=>X"00",
26899=>X"00",
26900=>X"00",
26901=>X"00",
26902=>X"00",
26903=>X"00",
26904=>X"00",
26905=>X"00",
26906=>X"00",
26907=>X"00",
26908=>X"00",
26909=>X"00",
26910=>X"00",
26911=>X"00",
26912=>X"00",
26913=>X"00",
26914=>X"00",
26915=>X"00",
26916=>X"00",
26917=>X"00",
26918=>X"00",
26919=>X"00",
26920=>X"00",
26921=>X"00",
26922=>X"00",
26923=>X"00",
26924=>X"00",
26925=>X"00",
26926=>X"00",
26927=>X"00",
26928=>X"00",
26929=>X"00",
26930=>X"00",
26931=>X"00",
26932=>X"00",
26933=>X"00",
26934=>X"00",
26935=>X"00",
26936=>X"00",
26937=>X"00",
26938=>X"00",
26939=>X"00",
26940=>X"00",
26941=>X"00",
26942=>X"00",
26943=>X"00",
26944=>X"00",
26945=>X"00",
26946=>X"00",
26947=>X"00",
26948=>X"00",
26949=>X"00",
26950=>X"00",
26951=>X"00",
26952=>X"00",
26953=>X"00",
26954=>X"00",
26955=>X"00",
26956=>X"00",
26957=>X"00",
26958=>X"00",
26959=>X"00",
26960=>X"00",
26961=>X"00",
26962=>X"00",
26963=>X"00",
26964=>X"00",
26965=>X"00",
26966=>X"00",
26967=>X"00",
26968=>X"00",
26969=>X"00",
26970=>X"00",
26971=>X"00",
26972=>X"00",
26973=>X"00",
26974=>X"00",
26975=>X"00",
26976=>X"00",
26977=>X"00",
26978=>X"00",
26979=>X"00",
26980=>X"00",
26981=>X"00",
26982=>X"00",
26983=>X"00",
26984=>X"00",
26985=>X"00",
26986=>X"00",
26987=>X"00",
26988=>X"00",
26989=>X"00",
26990=>X"00",
26991=>X"00",
26992=>X"00",
26993=>X"00",
26994=>X"00",
26995=>X"00",
26996=>X"00",
26997=>X"00",
26998=>X"00",
26999=>X"00",
27000=>X"00",
27001=>X"00",
27002=>X"00",
27003=>X"00",
27004=>X"00",
27005=>X"00",
27006=>X"00",
27007=>X"00",
27008=>X"00",
27009=>X"00",
27010=>X"00",
27011=>X"00",
27012=>X"00",
27013=>X"00",
27014=>X"00",
27015=>X"00",
27016=>X"00",
27017=>X"00",
27018=>X"00",
27019=>X"00",
27020=>X"00",
27021=>X"00",
27022=>X"00",
27023=>X"00",
27024=>X"00",
27025=>X"00",
27026=>X"00",
27027=>X"00",
27028=>X"00",
27029=>X"00",
27030=>X"00",
27031=>X"00",
27032=>X"00",
27033=>X"00",
27034=>X"00",
27035=>X"00",
27036=>X"00",
27037=>X"00",
27038=>X"00",
27039=>X"00",
27040=>X"00",
27041=>X"00",
27042=>X"00",
27043=>X"00",
27044=>X"00",
27045=>X"00",
27046=>X"00",
27047=>X"00",
27048=>X"00",
27049=>X"00",
27050=>X"00",
27051=>X"00",
27052=>X"00",
27053=>X"00",
27054=>X"00",
27055=>X"00",
27056=>X"00",
27057=>X"00",
27058=>X"00",
27059=>X"00",
27060=>X"00",
27061=>X"00",
27062=>X"00",
27063=>X"00",
27064=>X"00",
27065=>X"00",
27066=>X"00",
27067=>X"00",
27068=>X"00",
27069=>X"00",
27070=>X"00",
27071=>X"00",
27072=>X"00",
27073=>X"00",
27074=>X"00",
27075=>X"00",
27076=>X"00",
27077=>X"00",
27078=>X"00",
27079=>X"00",
27080=>X"00",
27081=>X"00",
27082=>X"00",
27083=>X"00",
27084=>X"00",
27085=>X"00",
27086=>X"00",
27087=>X"00",
27088=>X"00",
27089=>X"00",
27090=>X"00",
27091=>X"00",
27092=>X"00",
27093=>X"00",
27094=>X"00",
27095=>X"00",
27096=>X"00",
27097=>X"00",
27098=>X"00",
27099=>X"00",
27100=>X"00",
27101=>X"00",
27102=>X"00",
27103=>X"00",
27104=>X"00",
27105=>X"00",
27106=>X"00",
27107=>X"00",
27108=>X"00",
27109=>X"00",
27110=>X"00",
27111=>X"00",
27112=>X"00",
27113=>X"00",
27114=>X"00",
27115=>X"00",
27116=>X"00",
27117=>X"00",
27118=>X"00",
27119=>X"00",
27120=>X"00",
27121=>X"00",
27122=>X"00",
27123=>X"00",
27124=>X"00",
27125=>X"00",
27126=>X"00",
27127=>X"00",
27128=>X"00",
27129=>X"00",
27130=>X"00",
27131=>X"00",
27132=>X"00",
27133=>X"00",
27134=>X"00",
27135=>X"00",
27136=>X"00",
27137=>X"00",
27138=>X"00",
27139=>X"00",
27140=>X"00",
27141=>X"00",
27142=>X"00",
27143=>X"00",
27144=>X"00",
27145=>X"00",
27146=>X"00",
27147=>X"00",
27148=>X"00",
27149=>X"00",
27150=>X"00",
27151=>X"00",
27152=>X"00",
27153=>X"00",
27154=>X"00",
27155=>X"00",
27156=>X"00",
27157=>X"00",
27158=>X"00",
27159=>X"00",
27160=>X"00",
27161=>X"00",
27162=>X"00",
27163=>X"00",
27164=>X"00",
27165=>X"00",
27166=>X"00",
27167=>X"00",
27168=>X"00",
27169=>X"00",
27170=>X"00",
27171=>X"00",
27172=>X"00",
27173=>X"00",
27174=>X"00",
27175=>X"00",
27176=>X"00",
27177=>X"00",
27178=>X"00",
27179=>X"00",
27180=>X"00",
27181=>X"00",
27182=>X"00",
27183=>X"00",
27184=>X"00",
27185=>X"00",
27186=>X"00",
27187=>X"00",
27188=>X"00",
27189=>X"00",
27190=>X"00",
27191=>X"00",
27192=>X"00",
27193=>X"00",
27194=>X"00",
27195=>X"00",
27196=>X"00",
27197=>X"00",
27198=>X"00",
27199=>X"00",
27200=>X"00",
27201=>X"00",
27202=>X"00",
27203=>X"00",
27204=>X"00",
27205=>X"00",
27206=>X"00",
27207=>X"00",
27208=>X"00",
27209=>X"00",
27210=>X"00",
27211=>X"00",
27212=>X"00",
27213=>X"00",
27214=>X"00",
27215=>X"00",
27216=>X"00",
27217=>X"00",
27218=>X"00",
27219=>X"00",
27220=>X"00",
27221=>X"00",
27222=>X"00",
27223=>X"00",
27224=>X"00",
27225=>X"00",
27226=>X"00",
27227=>X"00",
27228=>X"00",
27229=>X"00",
27230=>X"00",
27231=>X"00",
27232=>X"00",
27233=>X"00",
27234=>X"00",
27235=>X"00",
27236=>X"00",
27237=>X"00",
27238=>X"00",
27239=>X"00",
27240=>X"00",
27241=>X"00",
27242=>X"00",
27243=>X"00",
27244=>X"00",
27245=>X"00",
27246=>X"00",
27247=>X"00",
27248=>X"00",
27249=>X"00",
27250=>X"00",
27251=>X"00",
27252=>X"00",
27253=>X"00",
27254=>X"00",
27255=>X"00",
27256=>X"00",
27257=>X"00",
27258=>X"00",
27259=>X"00",
27260=>X"00",
27261=>X"00",
27262=>X"00",
27263=>X"00",
27264=>X"00",
27265=>X"00",
27266=>X"00",
27267=>X"00",
27268=>X"00",
27269=>X"00",
27270=>X"00",
27271=>X"00",
27272=>X"00",
27273=>X"00",
27274=>X"00",
27275=>X"00",
27276=>X"00",
27277=>X"00",
27278=>X"00",
27279=>X"00",
27280=>X"00",
27281=>X"00",
27282=>X"00",
27283=>X"00",
27284=>X"00",
27285=>X"00",
27286=>X"00",
27287=>X"00",
27288=>X"00",
27289=>X"00",
27290=>X"00",
27291=>X"00",
27292=>X"00",
27293=>X"00",
27294=>X"00",
27295=>X"00",
27296=>X"00",
27297=>X"00",
27298=>X"00",
27299=>X"00",
27300=>X"00",
27301=>X"00",
27302=>X"00",
27303=>X"00",
27304=>X"00",
27305=>X"00",
27306=>X"00",
27307=>X"00",
27308=>X"00",
27309=>X"00",
27310=>X"00",
27311=>X"00",
27312=>X"00",
27313=>X"00",
27314=>X"00",
27315=>X"00",
27316=>X"00",
27317=>X"00",
27318=>X"00",
27319=>X"00",
27320=>X"00",
27321=>X"00",
27322=>X"00",
27323=>X"00",
27324=>X"00",
27325=>X"00",
27326=>X"00",
27327=>X"00",
27328=>X"00",
27329=>X"00",
27330=>X"00",
27331=>X"00",
27332=>X"00",
27333=>X"00",
27334=>X"00",
27335=>X"00",
27336=>X"00",
27337=>X"00",
27338=>X"00",
27339=>X"00",
27340=>X"00",
27341=>X"00",
27342=>X"00",
27343=>X"00",
27344=>X"00",
27345=>X"00",
27346=>X"00",
27347=>X"00",
27348=>X"00",
27349=>X"00",
27350=>X"00",
27351=>X"00",
27352=>X"00",
27353=>X"00",
27354=>X"00",
27355=>X"00",
27356=>X"00",
27357=>X"00",
27358=>X"00",
27359=>X"00",
27360=>X"00",
27361=>X"00",
27362=>X"00",
27363=>X"00",
27364=>X"00",
27365=>X"00",
27366=>X"00",
27367=>X"00",
27368=>X"00",
27369=>X"00",
27370=>X"00",
27371=>X"00",
27372=>X"00",
27373=>X"00",
27374=>X"00",
27375=>X"00",
27376=>X"00",
27377=>X"00",
27378=>X"00",
27379=>X"00",
27380=>X"00",
27381=>X"00",
27382=>X"00",
27383=>X"00",
27384=>X"00",
27385=>X"00",
27386=>X"00",
27387=>X"00",
27388=>X"00",
27389=>X"00",
27390=>X"00",
27391=>X"00",
27392=>X"00",
27393=>X"00",
27394=>X"00",
27395=>X"00",
27396=>X"00",
27397=>X"00",
27398=>X"00",
27399=>X"00",
27400=>X"00",
27401=>X"00",
27402=>X"00",
27403=>X"00",
27404=>X"00",
27405=>X"00",
27406=>X"00",
27407=>X"00",
27408=>X"00",
27409=>X"00",
27410=>X"00",
27411=>X"00",
27412=>X"00",
27413=>X"00",
27414=>X"00",
27415=>X"00",
27416=>X"00",
27417=>X"00",
27418=>X"00",
27419=>X"00",
27420=>X"00",
27421=>X"00",
27422=>X"00",
27423=>X"00",
27424=>X"00",
27425=>X"00",
27426=>X"00",
27427=>X"00",
27428=>X"00",
27429=>X"00",
27430=>X"00",
27431=>X"00",
27432=>X"00",
27433=>X"00",
27434=>X"00",
27435=>X"00",
27436=>X"00",
27437=>X"00",
27438=>X"00",
27439=>X"00",
27440=>X"00",
27441=>X"00",
27442=>X"00",
27443=>X"00",
27444=>X"00",
27445=>X"00",
27446=>X"00",
27447=>X"00",
27448=>X"00",
27449=>X"00",
27450=>X"00",
27451=>X"00",
27452=>X"00",
27453=>X"00",
27454=>X"00",
27455=>X"00",
27456=>X"00",
27457=>X"00",
27458=>X"00",
27459=>X"00",
27460=>X"00",
27461=>X"00",
27462=>X"00",
27463=>X"00",
27464=>X"00",
27465=>X"00",
27466=>X"00",
27467=>X"00",
27468=>X"00",
27469=>X"00",
27470=>X"00",
27471=>X"00",
27472=>X"00",
27473=>X"00",
27474=>X"00",
27475=>X"00",
27476=>X"00",
27477=>X"00",
27478=>X"00",
27479=>X"00",
27480=>X"00",
27481=>X"00",
27482=>X"00",
27483=>X"00",
27484=>X"00",
27485=>X"00",
27486=>X"00",
27487=>X"00",
27488=>X"00",
27489=>X"00",
27490=>X"00",
27491=>X"00",
27492=>X"00",
27493=>X"00",
27494=>X"00",
27495=>X"00",
27496=>X"00",
27497=>X"00",
27498=>X"00",
27499=>X"00",
27500=>X"00",
27501=>X"00",
27502=>X"00",
27503=>X"00",
27504=>X"00",
27505=>X"00",
27506=>X"00",
27507=>X"00",
27508=>X"00",
27509=>X"00",
27510=>X"00",
27511=>X"00",
27512=>X"00",
27513=>X"00",
27514=>X"00",
27515=>X"00",
27516=>X"00",
27517=>X"00",
27518=>X"00",
27519=>X"00",
27520=>X"00",
27521=>X"00",
27522=>X"00",
27523=>X"00",
27524=>X"00",
27525=>X"00",
27526=>X"00",
27527=>X"00",
27528=>X"00",
27529=>X"00",
27530=>X"00",
27531=>X"00",
27532=>X"00",
27533=>X"00",
27534=>X"00",
27535=>X"00",
27536=>X"00",
27537=>X"00",
27538=>X"00",
27539=>X"00",
27540=>X"00",
27541=>X"00",
27542=>X"00",
27543=>X"00",
27544=>X"00",
27545=>X"00",
27546=>X"00",
27547=>X"00",
27548=>X"00",
27549=>X"00",
27550=>X"00",
27551=>X"00",
27552=>X"00",
27553=>X"00",
27554=>X"00",
27555=>X"00",
27556=>X"00",
27557=>X"00",
27558=>X"00",
27559=>X"00",
27560=>X"00",
27561=>X"00",
27562=>X"00",
27563=>X"00",
27564=>X"00",
27565=>X"00",
27566=>X"00",
27567=>X"00",
27568=>X"00",
27569=>X"00",
27570=>X"00",
27571=>X"00",
27572=>X"00",
27573=>X"00",
27574=>X"00",
27575=>X"00",
27576=>X"00",
27577=>X"00",
27578=>X"00",
27579=>X"00",
27580=>X"00",
27581=>X"00",
27582=>X"00",
27583=>X"00",
27584=>X"00",
27585=>X"00",
27586=>X"00",
27587=>X"00",
27588=>X"00",
27589=>X"00",
27590=>X"00",
27591=>X"00",
27592=>X"00",
27593=>X"00",
27594=>X"00",
27595=>X"00",
27596=>X"00",
27597=>X"00",
27598=>X"00",
27599=>X"00",
27600=>X"00",
27601=>X"00",
27602=>X"00",
27603=>X"00",
27604=>X"00",
27605=>X"00",
27606=>X"00",
27607=>X"00",
27608=>X"00",
27609=>X"00",
27610=>X"00",
27611=>X"00",
27612=>X"00",
27613=>X"00",
27614=>X"00",
27615=>X"00",
27616=>X"00",
27617=>X"00",
27618=>X"00",
27619=>X"00",
27620=>X"00",
27621=>X"00",
27622=>X"00",
27623=>X"00",
27624=>X"00",
27625=>X"00",
27626=>X"00",
27627=>X"00",
27628=>X"00",
27629=>X"00",
27630=>X"00",
27631=>X"00",
27632=>X"00",
27633=>X"00",
27634=>X"00",
27635=>X"00",
27636=>X"00",
27637=>X"00",
27638=>X"00",
27639=>X"00",
27640=>X"00",
27641=>X"00",
27642=>X"00",
27643=>X"00",
27644=>X"00",
27645=>X"00",
27646=>X"00",
27647=>X"00",
27648=>X"00",
27649=>X"00",
27650=>X"00",
27651=>X"00",
27652=>X"00",
27653=>X"00",
27654=>X"00",
27655=>X"00",
27656=>X"00",
27657=>X"00",
27658=>X"00",
27659=>X"00",
27660=>X"00",
27661=>X"00",
27662=>X"00",
27663=>X"00",
27664=>X"00",
27665=>X"00",
27666=>X"00",
27667=>X"00",
27668=>X"00",
27669=>X"00",
27670=>X"00",
27671=>X"00",
27672=>X"00",
27673=>X"00",
27674=>X"00",
27675=>X"00",
27676=>X"00",
27677=>X"00",
27678=>X"00",
27679=>X"00",
27680=>X"00",
27681=>X"00",
27682=>X"00",
27683=>X"00",
27684=>X"00",
27685=>X"00",
27686=>X"00",
27687=>X"00",
27688=>X"00",
27689=>X"00",
27690=>X"00",
27691=>X"00",
27692=>X"00",
27693=>X"00",
27694=>X"00",
27695=>X"00",
27696=>X"00",
27697=>X"00",
27698=>X"00",
27699=>X"00",
27700=>X"00",
27701=>X"00",
27702=>X"00",
27703=>X"00",
27704=>X"00",
27705=>X"00",
27706=>X"00",
27707=>X"00",
27708=>X"00",
27709=>X"00",
27710=>X"00",
27711=>X"00",
27712=>X"00",
27713=>X"00",
27714=>X"00",
27715=>X"00",
27716=>X"00",
27717=>X"00",
27718=>X"00",
27719=>X"00",
27720=>X"00",
27721=>X"00",
27722=>X"00",
27723=>X"00",
27724=>X"00",
27725=>X"00",
27726=>X"00",
27727=>X"00",
27728=>X"00",
27729=>X"00",
27730=>X"00",
27731=>X"00",
27732=>X"00",
27733=>X"00",
27734=>X"00",
27735=>X"00",
27736=>X"00",
27737=>X"00",
27738=>X"00",
27739=>X"00",
27740=>X"00",
27741=>X"00",
27742=>X"00",
27743=>X"00",
27744=>X"00",
27745=>X"00",
27746=>X"00",
27747=>X"00",
27748=>X"00",
27749=>X"00",
27750=>X"00",
27751=>X"00",
27752=>X"00",
27753=>X"00",
27754=>X"00",
27755=>X"00",
27756=>X"00",
27757=>X"00",
27758=>X"00",
27759=>X"00",
27760=>X"00",
27761=>X"00",
27762=>X"00",
27763=>X"00",
27764=>X"00",
27765=>X"00",
27766=>X"00",
27767=>X"00",
27768=>X"00",
27769=>X"00",
27770=>X"00",
27771=>X"00",
27772=>X"00",
27773=>X"00",
27774=>X"00",
27775=>X"00",
27776=>X"00",
27777=>X"00",
27778=>X"00",
27779=>X"00",
27780=>X"00",
27781=>X"00",
27782=>X"00",
27783=>X"00",
27784=>X"00",
27785=>X"00",
27786=>X"00",
27787=>X"00",
27788=>X"00",
27789=>X"00",
27790=>X"00",
27791=>X"00",
27792=>X"00",
27793=>X"00",
27794=>X"00",
27795=>X"00",
27796=>X"00",
27797=>X"00",
27798=>X"00",
27799=>X"00",
27800=>X"00",
27801=>X"00",
27802=>X"00",
27803=>X"00",
27804=>X"00",
27805=>X"00",
27806=>X"00",
27807=>X"00",
27808=>X"00",
27809=>X"00",
27810=>X"00",
27811=>X"00",
27812=>X"00",
27813=>X"00",
27814=>X"00",
27815=>X"00",
27816=>X"00",
27817=>X"00",
27818=>X"00",
27819=>X"00",
27820=>X"00",
27821=>X"00",
27822=>X"00",
27823=>X"00",
27824=>X"00",
27825=>X"00",
27826=>X"00",
27827=>X"00",
27828=>X"00",
27829=>X"00",
27830=>X"00",
27831=>X"00",
27832=>X"00",
27833=>X"00",
27834=>X"00",
27835=>X"00",
27836=>X"00",
27837=>X"00",
27838=>X"00",
27839=>X"00",
27840=>X"00",
27841=>X"00",
27842=>X"00",
27843=>X"00",
27844=>X"00",
27845=>X"00",
27846=>X"00",
27847=>X"00",
27848=>X"00",
27849=>X"00",
27850=>X"00",
27851=>X"00",
27852=>X"00",
27853=>X"00",
27854=>X"00",
27855=>X"00",
27856=>X"00",
27857=>X"00",
27858=>X"00",
27859=>X"00",
27860=>X"00",
27861=>X"00",
27862=>X"00",
27863=>X"00",
27864=>X"00",
27865=>X"00",
27866=>X"00",
27867=>X"00",
27868=>X"00",
27869=>X"00",
27870=>X"00",
27871=>X"00",
27872=>X"00",
27873=>X"00",
27874=>X"00",
27875=>X"00",
27876=>X"00",
27877=>X"00",
27878=>X"00",
27879=>X"00",
27880=>X"00",
27881=>X"00",
27882=>X"00",
27883=>X"00",
27884=>X"00",
27885=>X"00",
27886=>X"00",
27887=>X"00",
27888=>X"00",
27889=>X"00",
27890=>X"00",
27891=>X"00",
27892=>X"00",
27893=>X"00",
27894=>X"00",
27895=>X"00",
27896=>X"00",
27897=>X"00",
27898=>X"00",
27899=>X"00",
27900=>X"00",
27901=>X"00",
27902=>X"00",
27903=>X"00",
27904=>X"00",
27905=>X"00",
27906=>X"00",
27907=>X"00",
27908=>X"00",
27909=>X"00",
27910=>X"00",
27911=>X"00",
27912=>X"00",
27913=>X"00",
27914=>X"00",
27915=>X"00",
27916=>X"00",
27917=>X"00",
27918=>X"00",
27919=>X"00",
27920=>X"00",
27921=>X"00",
27922=>X"00",
27923=>X"00",
27924=>X"00",
27925=>X"00",
27926=>X"00",
27927=>X"00",
27928=>X"00",
27929=>X"00",
27930=>X"00",
27931=>X"00",
27932=>X"00",
27933=>X"00",
27934=>X"00",
27935=>X"00",
27936=>X"00",
27937=>X"00",
27938=>X"00",
27939=>X"00",
27940=>X"00",
27941=>X"00",
27942=>X"00",
27943=>X"00",
27944=>X"00",
27945=>X"00",
27946=>X"00",
27947=>X"00",
27948=>X"00",
27949=>X"00",
27950=>X"00",
27951=>X"00",
27952=>X"00",
27953=>X"00",
27954=>X"00",
27955=>X"00",
27956=>X"00",
27957=>X"00",
27958=>X"00",
27959=>X"00",
27960=>X"00",
27961=>X"00",
27962=>X"00",
27963=>X"00",
27964=>X"00",
27965=>X"00",
27966=>X"00",
27967=>X"00",
27968=>X"00",
27969=>X"00",
27970=>X"00",
27971=>X"00",
27972=>X"00",
27973=>X"00",
27974=>X"00",
27975=>X"00",
27976=>X"00",
27977=>X"00",
27978=>X"00",
27979=>X"00",
27980=>X"00",
27981=>X"00",
27982=>X"00",
27983=>X"00",
27984=>X"00",
27985=>X"00",
27986=>X"00",
27987=>X"00",
27988=>X"00",
27989=>X"00",
27990=>X"00",
27991=>X"00",
27992=>X"00",
27993=>X"00",
27994=>X"00",
27995=>X"00",
27996=>X"00",
27997=>X"00",
27998=>X"00",
27999=>X"00",
28000=>X"00",
28001=>X"00",
28002=>X"00",
28003=>X"00",
28004=>X"00",
28005=>X"00",
28006=>X"00",
28007=>X"00",
28008=>X"00",
28009=>X"00",
28010=>X"00",
28011=>X"00",
28012=>X"00",
28013=>X"00",
28014=>X"00",
28015=>X"00",
28016=>X"00",
28017=>X"00",
28018=>X"00",
28019=>X"00",
28020=>X"00",
28021=>X"00",
28022=>X"00",
28023=>X"00",
28024=>X"00",
28025=>X"00",
28026=>X"00",
28027=>X"00",
28028=>X"00",
28029=>X"00",
28030=>X"00",
28031=>X"00",
28032=>X"00",
28033=>X"00",
28034=>X"00",
28035=>X"00",
28036=>X"00",
28037=>X"00",
28038=>X"00",
28039=>X"00",
28040=>X"00",
28041=>X"00",
28042=>X"00",
28043=>X"00",
28044=>X"00",
28045=>X"00",
28046=>X"00",
28047=>X"00",
28048=>X"00",
28049=>X"00",
28050=>X"00",
28051=>X"00",
28052=>X"00",
28053=>X"00",
28054=>X"00",
28055=>X"00",
28056=>X"00",
28057=>X"00",
28058=>X"00",
28059=>X"00",
28060=>X"00",
28061=>X"00",
28062=>X"00",
28063=>X"00",
28064=>X"00",
28065=>X"00",
28066=>X"00",
28067=>X"00",
28068=>X"00",
28069=>X"00",
28070=>X"00",
28071=>X"00",
28072=>X"00",
28073=>X"00",
28074=>X"00",
28075=>X"00",
28076=>X"00",
28077=>X"00",
28078=>X"00",
28079=>X"00",
28080=>X"00",
28081=>X"00",
28082=>X"00",
28083=>X"00",
28084=>X"00",
28085=>X"00",
28086=>X"00",
28087=>X"00",
28088=>X"00",
28089=>X"00",
28090=>X"00",
28091=>X"00",
28092=>X"00",
28093=>X"00",
28094=>X"00",
28095=>X"00",
28096=>X"00",
28097=>X"00",
28098=>X"00",
28099=>X"00",
28100=>X"00",
28101=>X"00",
28102=>X"00",
28103=>X"00",
28104=>X"00",
28105=>X"00",
28106=>X"00",
28107=>X"00",
28108=>X"00",
28109=>X"00",
28110=>X"00",
28111=>X"00",
28112=>X"00",
28113=>X"00",
28114=>X"00",
28115=>X"00",
28116=>X"00",
28117=>X"00",
28118=>X"00",
28119=>X"00",
28120=>X"00",
28121=>X"00",
28122=>X"00",
28123=>X"00",
28124=>X"00",
28125=>X"00",
28126=>X"00",
28127=>X"00",
28128=>X"00",
28129=>X"00",
28130=>X"00",
28131=>X"00",
28132=>X"00",
28133=>X"00",
28134=>X"00",
28135=>X"00",
28136=>X"00",
28137=>X"00",
28138=>X"00",
28139=>X"00",
28140=>X"00",
28141=>X"00",
28142=>X"00",
28143=>X"00",
28144=>X"00",
28145=>X"00",
28146=>X"00",
28147=>X"00",
28148=>X"00",
28149=>X"00",
28150=>X"00",
28151=>X"00",
28152=>X"00",
28153=>X"00",
28154=>X"00",
28155=>X"00",
28156=>X"00",
28157=>X"00",
28158=>X"00",
28159=>X"00",
28160=>X"00",
28161=>X"00",
28162=>X"00",
28163=>X"00",
28164=>X"00",
28165=>X"00",
28166=>X"00",
28167=>X"00",
28168=>X"00",
28169=>X"00",
28170=>X"00",
28171=>X"00",
28172=>X"00",
28173=>X"00",
28174=>X"00",
28175=>X"00",
28176=>X"00",
28177=>X"00",
28178=>X"00",
28179=>X"00",
28180=>X"00",
28181=>X"00",
28182=>X"00",
28183=>X"00",
28184=>X"00",
28185=>X"00",
28186=>X"00",
28187=>X"00",
28188=>X"00",
28189=>X"00",
28190=>X"00",
28191=>X"00",
28192=>X"00",
28193=>X"00",
28194=>X"00",
28195=>X"00",
28196=>X"00",
28197=>X"00",
28198=>X"00",
28199=>X"00",
28200=>X"00",
28201=>X"00",
28202=>X"00",
28203=>X"00",
28204=>X"00",
28205=>X"00",
28206=>X"00",
28207=>X"00",
28208=>X"00",
28209=>X"00",
28210=>X"00",
28211=>X"00",
28212=>X"00",
28213=>X"00",
28214=>X"00",
28215=>X"00",
28216=>X"00",
28217=>X"00",
28218=>X"00",
28219=>X"00",
28220=>X"00",
28221=>X"00",
28222=>X"00",
28223=>X"00",
28224=>X"00",
28225=>X"00",
28226=>X"00",
28227=>X"00",
28228=>X"00",
28229=>X"00",
28230=>X"00",
28231=>X"00",
28232=>X"00",
28233=>X"00",
28234=>X"00",
28235=>X"00",
28236=>X"00",
28237=>X"00",
28238=>X"00",
28239=>X"00",
28240=>X"00",
28241=>X"00",
28242=>X"00",
28243=>X"00",
28244=>X"00",
28245=>X"00",
28246=>X"00",
28247=>X"00",
28248=>X"00",
28249=>X"00",
28250=>X"00",
28251=>X"00",
28252=>X"00",
28253=>X"00",
28254=>X"00",
28255=>X"00",
28256=>X"00",
28257=>X"00",
28258=>X"00",
28259=>X"00",
28260=>X"00",
28261=>X"00",
28262=>X"00",
28263=>X"00",
28264=>X"00",
28265=>X"00",
28266=>X"00",
28267=>X"00",
28268=>X"00",
28269=>X"00",
28270=>X"00",
28271=>X"00",
28272=>X"00",
28273=>X"00",
28274=>X"00",
28275=>X"00",
28276=>X"00",
28277=>X"00",
28278=>X"00",
28279=>X"00",
28280=>X"00",
28281=>X"00",
28282=>X"00",
28283=>X"00",
28284=>X"00",
28285=>X"00",
28286=>X"00",
28287=>X"00",
28288=>X"00",
28289=>X"00",
28290=>X"00",
28291=>X"00",
28292=>X"00",
28293=>X"00",
28294=>X"00",
28295=>X"00",
28296=>X"00",
28297=>X"00",
28298=>X"00",
28299=>X"00",
28300=>X"00",
28301=>X"00",
28302=>X"00",
28303=>X"00",
28304=>X"00",
28305=>X"00",
28306=>X"00",
28307=>X"00",
28308=>X"00",
28309=>X"00",
28310=>X"00",
28311=>X"00",
28312=>X"00",
28313=>X"00",
28314=>X"00",
28315=>X"00",
28316=>X"00",
28317=>X"00",
28318=>X"00",
28319=>X"00",
28320=>X"00",
28321=>X"00",
28322=>X"00",
28323=>X"00",
28324=>X"00",
28325=>X"00",
28326=>X"00",
28327=>X"00",
28328=>X"00",
28329=>X"00",
28330=>X"00",
28331=>X"00",
28332=>X"00",
28333=>X"00",
28334=>X"00",
28335=>X"00",
28336=>X"00",
28337=>X"00",
28338=>X"00",
28339=>X"00",
28340=>X"00",
28341=>X"00",
28342=>X"00",
28343=>X"00",
28344=>X"00",
28345=>X"00",
28346=>X"00",
28347=>X"00",
28348=>X"00",
28349=>X"00",
28350=>X"00",
28351=>X"00",
28352=>X"00",
28353=>X"00",
28354=>X"00",
28355=>X"00",
28356=>X"00",
28357=>X"00",
28358=>X"00",
28359=>X"00",
28360=>X"00",
28361=>X"00",
28362=>X"00",
28363=>X"00",
28364=>X"00",
28365=>X"00",
28366=>X"00",
28367=>X"00",
28368=>X"00",
28369=>X"00",
28370=>X"00",
28371=>X"00",
28372=>X"00",
28373=>X"00",
28374=>X"00",
28375=>X"00",
28376=>X"00",
28377=>X"00",
28378=>X"00",
28379=>X"00",
28380=>X"00",
28381=>X"00",
28382=>X"00",
28383=>X"00",
28384=>X"00",
28385=>X"00",
28386=>X"00",
28387=>X"00",
28388=>X"00",
28389=>X"00",
28390=>X"00",
28391=>X"00",
28392=>X"00",
28393=>X"00",
28394=>X"00",
28395=>X"00",
28396=>X"00",
28397=>X"00",
28398=>X"00",
28399=>X"00",
28400=>X"00",
28401=>X"00",
28402=>X"00",
28403=>X"00",
28404=>X"00",
28405=>X"00",
28406=>X"00",
28407=>X"00",
28408=>X"00",
28409=>X"00",
28410=>X"00",
28411=>X"00",
28412=>X"00",
28413=>X"00",
28414=>X"00",
28415=>X"00",
28416=>X"00",
28417=>X"00",
28418=>X"00",
28419=>X"00",
28420=>X"00",
28421=>X"00",
28422=>X"00",
28423=>X"00",
28424=>X"00",
28425=>X"00",
28426=>X"00",
28427=>X"00",
28428=>X"00",
28429=>X"00",
28430=>X"00",
28431=>X"00",
28432=>X"00",
28433=>X"00",
28434=>X"00",
28435=>X"00",
28436=>X"00",
28437=>X"00",
28438=>X"00",
28439=>X"00",
28440=>X"00",
28441=>X"00",
28442=>X"00",
28443=>X"00",
28444=>X"00",
28445=>X"00",
28446=>X"00",
28447=>X"00",
28448=>X"00",
28449=>X"00",
28450=>X"00",
28451=>X"00",
28452=>X"00",
28453=>X"00",
28454=>X"00",
28455=>X"00",
28456=>X"00",
28457=>X"00",
28458=>X"00",
28459=>X"00",
28460=>X"00",
28461=>X"00",
28462=>X"00",
28463=>X"00",
28464=>X"00",
28465=>X"00",
28466=>X"00",
28467=>X"00",
28468=>X"00",
28469=>X"00",
28470=>X"00",
28471=>X"00",
28472=>X"00",
28473=>X"00",
28474=>X"00",
28475=>X"00",
28476=>X"00",
28477=>X"00",
28478=>X"00",
28479=>X"00",
28480=>X"00",
28481=>X"00",
28482=>X"00",
28483=>X"00",
28484=>X"00",
28485=>X"00",
28486=>X"00",
28487=>X"00",
28488=>X"00",
28489=>X"00",
28490=>X"00",
28491=>X"00",
28492=>X"00",
28493=>X"00",
28494=>X"00",
28495=>X"00",
28496=>X"00",
28497=>X"00",
28498=>X"00",
28499=>X"00",
28500=>X"00",
28501=>X"00",
28502=>X"00",
28503=>X"00",
28504=>X"00",
28505=>X"00",
28506=>X"00",
28507=>X"00",
28508=>X"00",
28509=>X"00",
28510=>X"00",
28511=>X"00",
28512=>X"00",
28513=>X"00",
28514=>X"00",
28515=>X"00",
28516=>X"00",
28517=>X"00",
28518=>X"00",
28519=>X"00",
28520=>X"00",
28521=>X"00",
28522=>X"00",
28523=>X"00",
28524=>X"00",
28525=>X"00",
28526=>X"00",
28527=>X"00",
28528=>X"00",
28529=>X"00",
28530=>X"00",
28531=>X"00",
28532=>X"00",
28533=>X"00",
28534=>X"00",
28535=>X"00",
28536=>X"00",
28537=>X"00",
28538=>X"00",
28539=>X"00",
28540=>X"00",
28541=>X"00",
28542=>X"00",
28543=>X"00",
28544=>X"00",
28545=>X"00",
28546=>X"00",
28547=>X"00",
28548=>X"00",
28549=>X"00",
28550=>X"00",
28551=>X"00",
28552=>X"00",
28553=>X"00",
28554=>X"00",
28555=>X"00",
28556=>X"00",
28557=>X"00",
28558=>X"00",
28559=>X"00",
28560=>X"00",
28561=>X"00",
28562=>X"00",
28563=>X"00",
28564=>X"00",
28565=>X"00",
28566=>X"00",
28567=>X"00",
28568=>X"00",
28569=>X"00",
28570=>X"00",
28571=>X"00",
28572=>X"00",
28573=>X"00",
28574=>X"00",
28575=>X"00",
28576=>X"00",
28577=>X"00",
28578=>X"00",
28579=>X"00",
28580=>X"00",
28581=>X"00",
28582=>X"00",
28583=>X"00",
28584=>X"00",
28585=>X"00",
28586=>X"00",
28587=>X"00",
28588=>X"00",
28589=>X"00",
28590=>X"00",
28591=>X"00",
28592=>X"00",
28593=>X"00",
28594=>X"00",
28595=>X"00",
28596=>X"00",
28597=>X"00",
28598=>X"00",
28599=>X"00",
28600=>X"00",
28601=>X"00",
28602=>X"00",
28603=>X"00",
28604=>X"00",
28605=>X"00",
28606=>X"00",
28607=>X"00",
28608=>X"00",
28609=>X"00",
28610=>X"00",
28611=>X"00",
28612=>X"00",
28613=>X"00",
28614=>X"00",
28615=>X"00",
28616=>X"00",
28617=>X"00",
28618=>X"00",
28619=>X"00",
28620=>X"00",
28621=>X"00",
28622=>X"00",
28623=>X"00",
28624=>X"00",
28625=>X"00",
28626=>X"00",
28627=>X"00",
28628=>X"00",
28629=>X"00",
28630=>X"00",
28631=>X"00",
28632=>X"00",
28633=>X"00",
28634=>X"00",
28635=>X"00",
28636=>X"00",
28637=>X"00",
28638=>X"00",
28639=>X"00",
28640=>X"00",
28641=>X"00",
28642=>X"00",
28643=>X"00",
28644=>X"00",
28645=>X"00",
28646=>X"00",
28647=>X"00",
28648=>X"00",
28649=>X"00",
28650=>X"00",
28651=>X"00",
28652=>X"00",
28653=>X"00",
28654=>X"00",
28655=>X"00",
28656=>X"00",
28657=>X"00",
28658=>X"00",
28659=>X"00",
28660=>X"00",
28661=>X"00",
28662=>X"00",
28663=>X"00",
28664=>X"00",
28665=>X"00",
28666=>X"00",
28667=>X"00",
28668=>X"00",
28669=>X"00",
28670=>X"00",
28671=>X"00",
28672=>X"00",
28673=>X"00",
28674=>X"00",
28675=>X"00",
28676=>X"00",
28677=>X"00",
28678=>X"00",
28679=>X"00",
28680=>X"00",
28681=>X"00",
28682=>X"00",
28683=>X"00",
28684=>X"00",
28685=>X"00",
28686=>X"00",
28687=>X"00",
28688=>X"00",
28689=>X"00",
28690=>X"00",
28691=>X"00",
28692=>X"00",
28693=>X"00",
28694=>X"00",
28695=>X"00",
28696=>X"00",
28697=>X"00",
28698=>X"00",
28699=>X"00",
28700=>X"00",
28701=>X"00",
28702=>X"00",
28703=>X"00",
28704=>X"00",
28705=>X"00",
28706=>X"00",
28707=>X"00",
28708=>X"00",
28709=>X"00",
28710=>X"00",
28711=>X"00",
28712=>X"00",
28713=>X"00",
28714=>X"00",
28715=>X"00",
28716=>X"00",
28717=>X"00",
28718=>X"00",
28719=>X"00",
28720=>X"00",
28721=>X"00",
28722=>X"00",
28723=>X"00",
28724=>X"00",
28725=>X"00",
28726=>X"00",
28727=>X"00",
28728=>X"00",
28729=>X"00",
28730=>X"00",
28731=>X"00",
28732=>X"00",
28733=>X"00",
28734=>X"00",
28735=>X"00",
28736=>X"00",
28737=>X"00",
28738=>X"00",
28739=>X"00",
28740=>X"00",
28741=>X"00",
28742=>X"00",
28743=>X"00",
28744=>X"00",
28745=>X"00",
28746=>X"00",
28747=>X"00",
28748=>X"00",
28749=>X"00",
28750=>X"00",
28751=>X"00",
28752=>X"00",
28753=>X"00",
28754=>X"00",
28755=>X"00",
28756=>X"00",
28757=>X"00",
28758=>X"00",
28759=>X"00",
28760=>X"00",
28761=>X"00",
28762=>X"00",
28763=>X"00",
28764=>X"00",
28765=>X"00",
28766=>X"00",
28767=>X"00",
28768=>X"00",
28769=>X"00",
28770=>X"00",
28771=>X"00",
28772=>X"00",
28773=>X"00",
28774=>X"00",
28775=>X"00",
28776=>X"00",
28777=>X"00",
28778=>X"00",
28779=>X"00",
28780=>X"00",
28781=>X"00",
28782=>X"00",
28783=>X"00",
28784=>X"00",
28785=>X"00",
28786=>X"00",
28787=>X"00",
28788=>X"00",
28789=>X"00",
28790=>X"00",
28791=>X"00",
28792=>X"00",
28793=>X"00",
28794=>X"00",
28795=>X"00",
28796=>X"00",
28797=>X"00",
28798=>X"00",
28799=>X"00",
28800=>X"00",
28801=>X"00",
28802=>X"00",
28803=>X"00",
28804=>X"00",
28805=>X"00",
28806=>X"00",
28807=>X"00",
28808=>X"00",
28809=>X"00",
28810=>X"00",
28811=>X"00",
28812=>X"00",
28813=>X"00",
28814=>X"00",
28815=>X"00",
28816=>X"00",
28817=>X"00",
28818=>X"00",
28819=>X"00",
28820=>X"00",
28821=>X"00",
28822=>X"00",
28823=>X"00",
28824=>X"00",
28825=>X"00",
28826=>X"00",
28827=>X"00",
28828=>X"00",
28829=>X"00",
28830=>X"00",
28831=>X"00",
28832=>X"00",
28833=>X"00",
28834=>X"00",
28835=>X"00",
28836=>X"00",
28837=>X"00",
28838=>X"00",
28839=>X"00",
28840=>X"00",
28841=>X"00",
28842=>X"00",
28843=>X"00",
28844=>X"00",
28845=>X"00",
28846=>X"00",
28847=>X"00",
28848=>X"00",
28849=>X"00",
28850=>X"00",
28851=>X"00",
28852=>X"00",
28853=>X"00",
28854=>X"00",
28855=>X"00",
28856=>X"00",
28857=>X"00",
28858=>X"00",
28859=>X"00",
28860=>X"00",
28861=>X"00",
28862=>X"00",
28863=>X"00",
28864=>X"00",
28865=>X"00",
28866=>X"00",
28867=>X"00",
28868=>X"00",
28869=>X"00",
28870=>X"00",
28871=>X"00",
28872=>X"00",
28873=>X"00",
28874=>X"00",
28875=>X"00",
28876=>X"00",
28877=>X"00",
28878=>X"00",
28879=>X"00",
28880=>X"00",
28881=>X"00",
28882=>X"00",
28883=>X"00",
28884=>X"00",
28885=>X"00",
28886=>X"00",
28887=>X"00",
28888=>X"00",
28889=>X"00",
28890=>X"00",
28891=>X"00",
28892=>X"00",
28893=>X"00",
28894=>X"00",
28895=>X"00",
28896=>X"00",
28897=>X"00",
28898=>X"00",
28899=>X"00",
28900=>X"00",
28901=>X"00",
28902=>X"00",
28903=>X"00",
28904=>X"00",
28905=>X"00",
28906=>X"00",
28907=>X"00",
28908=>X"00",
28909=>X"00",
28910=>X"00",
28911=>X"00",
28912=>X"00",
28913=>X"00",
28914=>X"00",
28915=>X"00",
28916=>X"00",
28917=>X"00",
28918=>X"00",
28919=>X"00",
28920=>X"00",
28921=>X"00",
28922=>X"00",
28923=>X"00",
28924=>X"00",
28925=>X"00",
28926=>X"00",
28927=>X"00",
28928=>X"00",
28929=>X"00",
28930=>X"00",
28931=>X"00",
28932=>X"00",
28933=>X"00",
28934=>X"00",
28935=>X"00",
28936=>X"00",
28937=>X"00",
28938=>X"00",
28939=>X"00",
28940=>X"00",
28941=>X"00",
28942=>X"00",
28943=>X"00",
28944=>X"00",
28945=>X"00",
28946=>X"00",
28947=>X"00",
28948=>X"00",
28949=>X"00",
28950=>X"00",
28951=>X"00",
28952=>X"00",
28953=>X"00",
28954=>X"00",
28955=>X"00",
28956=>X"00",
28957=>X"00",
28958=>X"00",
28959=>X"00",
28960=>X"00",
28961=>X"00",
28962=>X"00",
28963=>X"00",
28964=>X"00",
28965=>X"00",
28966=>X"00",
28967=>X"00",
28968=>X"00",
28969=>X"00",
28970=>X"00",
28971=>X"00",
28972=>X"00",
28973=>X"00",
28974=>X"00",
28975=>X"00",
28976=>X"00",
28977=>X"00",
28978=>X"00",
28979=>X"00",
28980=>X"00",
28981=>X"00",
28982=>X"00",
28983=>X"00",
28984=>X"00",
28985=>X"00",
28986=>X"00",
28987=>X"00",
28988=>X"00",
28989=>X"00",
28990=>X"00",
28991=>X"00",
28992=>X"00",
28993=>X"00",
28994=>X"00",
28995=>X"00",
28996=>X"00",
28997=>X"00",
28998=>X"00",
28999=>X"00",
29000=>X"00",
29001=>X"00",
29002=>X"00",
29003=>X"00",
29004=>X"00",
29005=>X"00",
29006=>X"00",
29007=>X"00",
29008=>X"00",
29009=>X"00",
29010=>X"00",
29011=>X"00",
29012=>X"00",
29013=>X"00",
29014=>X"00",
29015=>X"00",
29016=>X"00",
29017=>X"00",
29018=>X"00",
29019=>X"00",
29020=>X"00",
29021=>X"00",
29022=>X"00",
29023=>X"00",
29024=>X"00",
29025=>X"00",
29026=>X"00",
29027=>X"00",
29028=>X"00",
29029=>X"00",
29030=>X"00",
29031=>X"00",
29032=>X"00",
29033=>X"00",
29034=>X"00",
29035=>X"00",
29036=>X"00",
29037=>X"00",
29038=>X"00",
29039=>X"00",
29040=>X"00",
29041=>X"00",
29042=>X"00",
29043=>X"00",
29044=>X"00",
29045=>X"00",
29046=>X"00",
29047=>X"00",
29048=>X"00",
29049=>X"00",
29050=>X"00",
29051=>X"00",
29052=>X"00",
29053=>X"00",
29054=>X"00",
29055=>X"00",
29056=>X"00",
29057=>X"00",
29058=>X"00",
29059=>X"00",
29060=>X"00",
29061=>X"00",
29062=>X"00",
29063=>X"00",
29064=>X"00",
29065=>X"00",
29066=>X"00",
29067=>X"00",
29068=>X"00",
29069=>X"00",
29070=>X"00",
29071=>X"00",
29072=>X"00",
29073=>X"00",
29074=>X"00",
29075=>X"00",
29076=>X"00",
29077=>X"00",
29078=>X"00",
29079=>X"00",
29080=>X"00",
29081=>X"00",
29082=>X"00",
29083=>X"00",
29084=>X"00",
29085=>X"00",
29086=>X"00",
29087=>X"00",
29088=>X"00",
29089=>X"00",
29090=>X"00",
29091=>X"00",
29092=>X"00",
29093=>X"00",
29094=>X"00",
29095=>X"00",
29096=>X"00",
29097=>X"00",
29098=>X"00",
29099=>X"00",
29100=>X"00",
29101=>X"00",
29102=>X"00",
29103=>X"00",
29104=>X"00",
29105=>X"00",
29106=>X"00",
29107=>X"00",
29108=>X"00",
29109=>X"00",
29110=>X"00",
29111=>X"00",
29112=>X"00",
29113=>X"00",
29114=>X"00",
29115=>X"00",
29116=>X"00",
29117=>X"00",
29118=>X"00",
29119=>X"00",
29120=>X"00",
29121=>X"00",
29122=>X"00",
29123=>X"00",
29124=>X"00",
29125=>X"00",
29126=>X"00",
29127=>X"00",
29128=>X"00",
29129=>X"00",
29130=>X"00",
29131=>X"00",
29132=>X"00",
29133=>X"00",
29134=>X"00",
29135=>X"00",
29136=>X"00",
29137=>X"00",
29138=>X"00",
29139=>X"00",
29140=>X"00",
29141=>X"00",
29142=>X"00",
29143=>X"00",
29144=>X"00",
29145=>X"00",
29146=>X"00",
29147=>X"00",
29148=>X"00",
29149=>X"00",
29150=>X"00",
29151=>X"00",
29152=>X"00",
29153=>X"00",
29154=>X"00",
29155=>X"00",
29156=>X"00",
29157=>X"00",
29158=>X"00",
29159=>X"00",
29160=>X"00",
29161=>X"00",
29162=>X"00",
29163=>X"00",
29164=>X"00",
29165=>X"00",
29166=>X"00",
29167=>X"00",
29168=>X"00",
29169=>X"00",
29170=>X"00",
29171=>X"00",
29172=>X"00",
29173=>X"00",
29174=>X"00",
29175=>X"00",
29176=>X"00",
29177=>X"00",
29178=>X"00",
29179=>X"00",
29180=>X"00",
29181=>X"00",
29182=>X"00",
29183=>X"00",
29184=>X"00",
29185=>X"00",
29186=>X"00",
29187=>X"00",
29188=>X"00",
29189=>X"00",
29190=>X"00",
29191=>X"00",
29192=>X"00",
29193=>X"00",
29194=>X"00",
29195=>X"00",
29196=>X"00",
29197=>X"00",
29198=>X"00",
29199=>X"00",
29200=>X"00",
29201=>X"00",
29202=>X"00",
29203=>X"00",
29204=>X"00",
29205=>X"00",
29206=>X"00",
29207=>X"00",
29208=>X"00",
29209=>X"00",
29210=>X"00",
29211=>X"00",
29212=>X"00",
29213=>X"00",
29214=>X"00",
29215=>X"00",
29216=>X"00",
29217=>X"00",
29218=>X"00",
29219=>X"00",
29220=>X"00",
29221=>X"00",
29222=>X"00",
29223=>X"00",
29224=>X"00",
29225=>X"00",
29226=>X"00",
29227=>X"00",
29228=>X"00",
29229=>X"00",
29230=>X"00",
29231=>X"00",
29232=>X"00",
29233=>X"00",
29234=>X"00",
29235=>X"00",
29236=>X"00",
29237=>X"00",
29238=>X"00",
29239=>X"00",
29240=>X"00",
29241=>X"00",
29242=>X"00",
29243=>X"00",
29244=>X"00",
29245=>X"00",
29246=>X"00",
29247=>X"00",
29248=>X"00",
29249=>X"00",
29250=>X"00",
29251=>X"00",
29252=>X"00",
29253=>X"00",
29254=>X"00",
29255=>X"00",
29256=>X"00",
29257=>X"00",
29258=>X"00",
29259=>X"00",
29260=>X"00",
29261=>X"00",
29262=>X"00",
29263=>X"00",
29264=>X"00",
29265=>X"00",
29266=>X"00",
29267=>X"00",
29268=>X"00",
29269=>X"00",
29270=>X"00",
29271=>X"00",
29272=>X"00",
29273=>X"00",
29274=>X"00",
29275=>X"00",
29276=>X"00",
29277=>X"00",
29278=>X"00",
29279=>X"00",
29280=>X"00",
29281=>X"00",
29282=>X"00",
29283=>X"00",
29284=>X"00",
29285=>X"00",
29286=>X"00",
29287=>X"00",
29288=>X"00",
29289=>X"00",
29290=>X"00",
29291=>X"00",
29292=>X"00",
29293=>X"00",
29294=>X"00",
29295=>X"00",
29296=>X"00",
29297=>X"00",
29298=>X"00",
29299=>X"00",
29300=>X"00",
29301=>X"00",
29302=>X"00",
29303=>X"00",
29304=>X"00",
29305=>X"00",
29306=>X"00",
29307=>X"00",
29308=>X"00",
29309=>X"00",
29310=>X"00",
29311=>X"00",
29312=>X"00",
29313=>X"00",
29314=>X"00",
29315=>X"00",
29316=>X"00",
29317=>X"00",
29318=>X"00",
29319=>X"00",
29320=>X"00",
29321=>X"00",
29322=>X"00",
29323=>X"00",
29324=>X"00",
29325=>X"00",
29326=>X"00",
29327=>X"00",
29328=>X"00",
29329=>X"00",
29330=>X"00",
29331=>X"00",
29332=>X"00",
29333=>X"00",
29334=>X"00",
29335=>X"00",
29336=>X"00",
29337=>X"00",
29338=>X"00",
29339=>X"00",
29340=>X"00",
29341=>X"00",
29342=>X"00",
29343=>X"00",
29344=>X"00",
29345=>X"00",
29346=>X"00",
29347=>X"00",
29348=>X"00",
29349=>X"00",
29350=>X"00",
29351=>X"00",
29352=>X"00",
29353=>X"00",
29354=>X"00",
29355=>X"00",
29356=>X"00",
29357=>X"00",
29358=>X"00",
29359=>X"00",
29360=>X"00",
29361=>X"00",
29362=>X"00",
29363=>X"00",
29364=>X"00",
29365=>X"00",
29366=>X"00",
29367=>X"00",
29368=>X"00",
29369=>X"00",
29370=>X"00",
29371=>X"00",
29372=>X"00",
29373=>X"00",
29374=>X"00",
29375=>X"00",
29376=>X"00",
29377=>X"00",
29378=>X"00",
29379=>X"00",
29380=>X"00",
29381=>X"00",
29382=>X"00",
29383=>X"00",
29384=>X"00",
29385=>X"00",
29386=>X"00",
29387=>X"00",
29388=>X"00",
29389=>X"00",
29390=>X"00",
29391=>X"00",
29392=>X"00",
29393=>X"00",
29394=>X"00",
29395=>X"00",
29396=>X"00",
29397=>X"00",
29398=>X"00",
29399=>X"00",
29400=>X"00",
29401=>X"00",
29402=>X"00",
29403=>X"00",
29404=>X"00",
29405=>X"00",
29406=>X"00",
29407=>X"00",
29408=>X"00",
29409=>X"00",
29410=>X"00",
29411=>X"00",
29412=>X"00",
29413=>X"00",
29414=>X"00",
29415=>X"00",
29416=>X"00",
29417=>X"00",
29418=>X"00",
29419=>X"00",
29420=>X"00",
29421=>X"00",
29422=>X"00",
29423=>X"00",
29424=>X"00",
29425=>X"00",
29426=>X"00",
29427=>X"00",
29428=>X"00",
29429=>X"00",
29430=>X"00",
29431=>X"00",
29432=>X"00",
29433=>X"00",
29434=>X"00",
29435=>X"00",
29436=>X"00",
29437=>X"00",
29438=>X"00",
29439=>X"00",
29440=>X"00",
29441=>X"00",
29442=>X"00",
29443=>X"00",
29444=>X"00",
29445=>X"00",
29446=>X"00",
29447=>X"00",
29448=>X"00",
29449=>X"00",
29450=>X"00",
29451=>X"00",
29452=>X"00",
29453=>X"00",
29454=>X"00",
29455=>X"00",
29456=>X"00",
29457=>X"00",
29458=>X"00",
29459=>X"00",
29460=>X"00",
29461=>X"00",
29462=>X"00",
29463=>X"00",
29464=>X"00",
29465=>X"00",
29466=>X"00",
29467=>X"00",
29468=>X"00",
29469=>X"00",
29470=>X"00",
29471=>X"00",
29472=>X"00",
29473=>X"00",
29474=>X"00",
29475=>X"00",
29476=>X"00",
29477=>X"00",
29478=>X"00",
29479=>X"00",
29480=>X"00",
29481=>X"00",
29482=>X"00",
29483=>X"00",
29484=>X"00",
29485=>X"00",
29486=>X"00",
29487=>X"00",
29488=>X"00",
29489=>X"00",
29490=>X"00",
29491=>X"00",
29492=>X"00",
29493=>X"00",
29494=>X"00",
29495=>X"00",
29496=>X"00",
29497=>X"00",
29498=>X"00",
29499=>X"00",
29500=>X"00",
29501=>X"00",
29502=>X"00",
29503=>X"00",
29504=>X"00",
29505=>X"00",
29506=>X"00",
29507=>X"00",
29508=>X"00",
29509=>X"00",
29510=>X"00",
29511=>X"00",
29512=>X"00",
29513=>X"00",
29514=>X"00",
29515=>X"00",
29516=>X"00",
29517=>X"00",
29518=>X"00",
29519=>X"00",
29520=>X"00",
29521=>X"00",
29522=>X"00",
29523=>X"00",
29524=>X"00",
29525=>X"00",
29526=>X"00",
29527=>X"00",
29528=>X"00",
29529=>X"00",
29530=>X"00",
29531=>X"00",
29532=>X"00",
29533=>X"00",
29534=>X"00",
29535=>X"00",
29536=>X"00",
29537=>X"00",
29538=>X"00",
29539=>X"00",
29540=>X"00",
29541=>X"00",
29542=>X"00",
29543=>X"00",
29544=>X"00",
29545=>X"00",
29546=>X"00",
29547=>X"00",
29548=>X"00",
29549=>X"00",
29550=>X"00",
29551=>X"00",
29552=>X"00",
29553=>X"00",
29554=>X"00",
29555=>X"00",
29556=>X"00",
29557=>X"00",
29558=>X"00",
29559=>X"00",
29560=>X"00",
29561=>X"00",
29562=>X"00",
29563=>X"00",
29564=>X"00",
29565=>X"00",
29566=>X"00",
29567=>X"00",
29568=>X"00",
29569=>X"00",
29570=>X"00",
29571=>X"00",
29572=>X"00",
29573=>X"00",
29574=>X"00",
29575=>X"00",
29576=>X"00",
29577=>X"00",
29578=>X"00",
29579=>X"00",
29580=>X"00",
29581=>X"00",
29582=>X"00",
29583=>X"00",
29584=>X"00",
29585=>X"00",
29586=>X"00",
29587=>X"00",
29588=>X"00",
29589=>X"00",
29590=>X"00",
29591=>X"00",
29592=>X"00",
29593=>X"00",
29594=>X"00",
29595=>X"00",
29596=>X"00",
29597=>X"00",
29598=>X"00",
29599=>X"00",
29600=>X"00",
29601=>X"00",
29602=>X"00",
29603=>X"00",
29604=>X"00",
29605=>X"00",
29606=>X"00",
29607=>X"00",
29608=>X"00",
29609=>X"00",
29610=>X"00",
29611=>X"00",
29612=>X"00",
29613=>X"00",
29614=>X"00",
29615=>X"00",
29616=>X"00",
29617=>X"00",
29618=>X"00",
29619=>X"00",
29620=>X"00",
29621=>X"00",
29622=>X"00",
29623=>X"00",
29624=>X"00",
29625=>X"00",
29626=>X"00",
29627=>X"00",
29628=>X"00",
29629=>X"00",
29630=>X"00",
29631=>X"00",
29632=>X"00",
29633=>X"00",
29634=>X"00",
29635=>X"00",
29636=>X"00",
29637=>X"00",
29638=>X"00",
29639=>X"00",
29640=>X"00",
29641=>X"00",
29642=>X"00",
29643=>X"00",
29644=>X"00",
29645=>X"00",
29646=>X"00",
29647=>X"00",
29648=>X"00",
29649=>X"00",
29650=>X"00",
29651=>X"00",
29652=>X"00",
29653=>X"00",
29654=>X"00",
29655=>X"00",
29656=>X"00",
29657=>X"00",
29658=>X"00",
29659=>X"00",
29660=>X"00",
29661=>X"00",
29662=>X"00",
29663=>X"00",
29664=>X"00",
29665=>X"00",
29666=>X"00",
29667=>X"00",
29668=>X"00",
29669=>X"00",
29670=>X"00",
29671=>X"00",
29672=>X"00",
29673=>X"00",
29674=>X"00",
29675=>X"00",
29676=>X"00",
29677=>X"00",
29678=>X"00",
29679=>X"00",
29680=>X"00",
29681=>X"00",
29682=>X"00",
29683=>X"00",
29684=>X"00",
29685=>X"00",
29686=>X"00",
29687=>X"00",
29688=>X"00",
29689=>X"00",
29690=>X"00",
29691=>X"00",
29692=>X"00",
29693=>X"00",
29694=>X"00",
29695=>X"00",
29696=>X"00",
29697=>X"00",
29698=>X"00",
29699=>X"00",
29700=>X"00",
29701=>X"00",
29702=>X"00",
29703=>X"00",
29704=>X"00",
29705=>X"00",
29706=>X"00",
29707=>X"00",
29708=>X"00",
29709=>X"00",
29710=>X"00",
29711=>X"00",
29712=>X"00",
29713=>X"00",
29714=>X"00",
29715=>X"00",
29716=>X"00",
29717=>X"00",
29718=>X"00",
29719=>X"00",
29720=>X"00",
29721=>X"00",
29722=>X"00",
29723=>X"00",
29724=>X"00",
29725=>X"00",
29726=>X"00",
29727=>X"00",
29728=>X"00",
29729=>X"00",
29730=>X"00",
29731=>X"00",
29732=>X"00",
29733=>X"00",
29734=>X"00",
29735=>X"00",
29736=>X"00",
29737=>X"00",
29738=>X"00",
29739=>X"00",
29740=>X"00",
29741=>X"00",
29742=>X"00",
29743=>X"00",
29744=>X"00",
29745=>X"00",
29746=>X"00",
29747=>X"00",
29748=>X"00",
29749=>X"00",
29750=>X"00",
29751=>X"00",
29752=>X"00",
29753=>X"00",
29754=>X"00",
29755=>X"00",
29756=>X"00",
29757=>X"00",
29758=>X"00",
29759=>X"00",
29760=>X"00",
29761=>X"00",
29762=>X"00",
29763=>X"00",
29764=>X"00",
29765=>X"00",
29766=>X"00",
29767=>X"00",
29768=>X"00",
29769=>X"00",
29770=>X"00",
29771=>X"00",
29772=>X"00",
29773=>X"00",
29774=>X"00",
29775=>X"00",
29776=>X"00",
29777=>X"00",
29778=>X"00",
29779=>X"00",
29780=>X"00",
29781=>X"00",
29782=>X"00",
29783=>X"00",
29784=>X"00",
29785=>X"00",
29786=>X"00",
29787=>X"00",
29788=>X"00",
29789=>X"00",
29790=>X"00",
29791=>X"00",
29792=>X"00",
29793=>X"00",
29794=>X"00",
29795=>X"00",
29796=>X"00",
29797=>X"00",
29798=>X"00",
29799=>X"00",
29800=>X"00",
29801=>X"00",
29802=>X"00",
29803=>X"00",
29804=>X"00",
29805=>X"00",
29806=>X"00",
29807=>X"00",
29808=>X"00",
29809=>X"00",
29810=>X"00",
29811=>X"00",
29812=>X"00",
29813=>X"00",
29814=>X"00",
29815=>X"00",
29816=>X"00",
29817=>X"00",
29818=>X"00",
29819=>X"00",
29820=>X"00",
29821=>X"00",
29822=>X"00",
29823=>X"00",
29824=>X"00",
29825=>X"00",
29826=>X"00",
29827=>X"00",
29828=>X"00",
29829=>X"00",
29830=>X"00",
29831=>X"00",
29832=>X"00",
29833=>X"00",
29834=>X"00",
29835=>X"00",
29836=>X"00",
29837=>X"00",
29838=>X"00",
29839=>X"00",
29840=>X"00",
29841=>X"00",
29842=>X"00",
29843=>X"00",
29844=>X"00",
29845=>X"00",
29846=>X"00",
29847=>X"00",
29848=>X"00",
29849=>X"00",
29850=>X"00",
29851=>X"00",
29852=>X"00",
29853=>X"00",
29854=>X"00",
29855=>X"00",
29856=>X"00",
29857=>X"00",
29858=>X"00",
29859=>X"00",
29860=>X"00",
29861=>X"00",
29862=>X"00",
29863=>X"00",
29864=>X"00",
29865=>X"00",
29866=>X"00",
29867=>X"00",
29868=>X"00",
29869=>X"00",
29870=>X"00",
29871=>X"00",
29872=>X"00",
29873=>X"00",
29874=>X"00",
29875=>X"00",
29876=>X"00",
29877=>X"00",
29878=>X"00",
29879=>X"00",
29880=>X"00",
29881=>X"00",
29882=>X"00",
29883=>X"00",
29884=>X"00",
29885=>X"00",
29886=>X"00",
29887=>X"00",
29888=>X"00",
29889=>X"00",
29890=>X"00",
29891=>X"00",
29892=>X"00",
29893=>X"00",
29894=>X"00",
29895=>X"00",
29896=>X"00",
29897=>X"00",
29898=>X"00",
29899=>X"00",
29900=>X"00",
29901=>X"00",
29902=>X"00",
29903=>X"00",
29904=>X"00",
29905=>X"00",
29906=>X"00",
29907=>X"00",
29908=>X"00",
29909=>X"00",
29910=>X"00",
29911=>X"00",
29912=>X"00",
29913=>X"00",
29914=>X"00",
29915=>X"00",
29916=>X"00",
29917=>X"00",
29918=>X"00",
29919=>X"00",
29920=>X"00",
29921=>X"00",
29922=>X"00",
29923=>X"00",
29924=>X"00",
29925=>X"00",
29926=>X"00",
29927=>X"00",
29928=>X"00",
29929=>X"00",
29930=>X"00",
29931=>X"00",
29932=>X"00",
29933=>X"00",
29934=>X"00",
29935=>X"00",
29936=>X"00",
29937=>X"00",
29938=>X"00",
29939=>X"00",
29940=>X"00",
29941=>X"00",
29942=>X"00",
29943=>X"00",
29944=>X"00",
29945=>X"00",
29946=>X"00",
29947=>X"00",
29948=>X"00",
29949=>X"00",
29950=>X"00",
29951=>X"00",
29952=>X"00",
29953=>X"00",
29954=>X"00",
29955=>X"00",
29956=>X"00",
29957=>X"00",
29958=>X"00",
29959=>X"00",
29960=>X"00",
29961=>X"00",
29962=>X"00",
29963=>X"00",
29964=>X"00",
29965=>X"00",
29966=>X"00",
29967=>X"00",
29968=>X"00",
29969=>X"00",
29970=>X"00",
29971=>X"00",
29972=>X"00",
29973=>X"00",
29974=>X"00",
29975=>X"00",
29976=>X"00",
29977=>X"00",
29978=>X"00",
29979=>X"00",
29980=>X"00",
29981=>X"00",
29982=>X"00",
29983=>X"00",
29984=>X"00",
29985=>X"00",
29986=>X"00",
29987=>X"00",
29988=>X"00",
29989=>X"00",
29990=>X"00",
29991=>X"00",
29992=>X"00",
29993=>X"00",
29994=>X"00",
29995=>X"00",
29996=>X"00",
29997=>X"00",
29998=>X"00",
29999=>X"00",
30000=>X"00",
30001=>X"00",
30002=>X"00",
30003=>X"00",
30004=>X"00",
30005=>X"00",
30006=>X"00",
30007=>X"00",
30008=>X"00",
30009=>X"00",
30010=>X"00",
30011=>X"00",
30012=>X"00",
30013=>X"00",
30014=>X"00",
30015=>X"00",
30016=>X"00",
30017=>X"00",
30018=>X"00",
30019=>X"00",
30020=>X"00",
30021=>X"00",
30022=>X"00",
30023=>X"00",
30024=>X"00",
30025=>X"00",
30026=>X"00",
30027=>X"00",
30028=>X"00",
30029=>X"00",
30030=>X"00",
30031=>X"00",
30032=>X"00",
30033=>X"00",
30034=>X"00",
30035=>X"00",
30036=>X"00",
30037=>X"00",
30038=>X"00",
30039=>X"00",
30040=>X"00",
30041=>X"00",
30042=>X"00",
30043=>X"00",
30044=>X"00",
30045=>X"00",
30046=>X"00",
30047=>X"00",
30048=>X"00",
30049=>X"00",
30050=>X"00",
30051=>X"00",
30052=>X"00",
30053=>X"00",
30054=>X"00",
30055=>X"00",
30056=>X"00",
30057=>X"00",
30058=>X"00",
30059=>X"00",
30060=>X"00",
30061=>X"00",
30062=>X"00",
30063=>X"00",
30064=>X"00",
30065=>X"00",
30066=>X"00",
30067=>X"00",
30068=>X"00",
30069=>X"00",
30070=>X"00",
30071=>X"00",
30072=>X"00",
30073=>X"00",
30074=>X"00",
30075=>X"00",
30076=>X"00",
30077=>X"00",
30078=>X"00",
30079=>X"00",
30080=>X"00",
30081=>X"00",
30082=>X"00",
30083=>X"00",
30084=>X"00",
30085=>X"00",
30086=>X"00",
30087=>X"00",
30088=>X"00",
30089=>X"00",
30090=>X"00",
30091=>X"00",
30092=>X"00",
30093=>X"00",
30094=>X"00",
30095=>X"00",
30096=>X"00",
30097=>X"00",
30098=>X"00",
30099=>X"00",
30100=>X"00",
30101=>X"00",
30102=>X"00",
30103=>X"00",
30104=>X"00",
30105=>X"00",
30106=>X"00",
30107=>X"00",
30108=>X"00",
30109=>X"00",
30110=>X"00",
30111=>X"00",
30112=>X"00",
30113=>X"00",
30114=>X"00",
30115=>X"00",
30116=>X"00",
30117=>X"00",
30118=>X"00",
30119=>X"00",
30120=>X"00",
30121=>X"00",
30122=>X"00",
30123=>X"00",
30124=>X"00",
30125=>X"00",
30126=>X"00",
30127=>X"00",
30128=>X"00",
30129=>X"00",
30130=>X"00",
30131=>X"00",
30132=>X"00",
30133=>X"00",
30134=>X"00",
30135=>X"00",
30136=>X"00",
30137=>X"00",
30138=>X"00",
30139=>X"00",
30140=>X"00",
30141=>X"00",
30142=>X"00",
30143=>X"00",
30144=>X"00",
30145=>X"00",
30146=>X"00",
30147=>X"00",
30148=>X"00",
30149=>X"00",
30150=>X"00",
30151=>X"00",
30152=>X"00",
30153=>X"00",
30154=>X"00",
30155=>X"00",
30156=>X"00",
30157=>X"00",
30158=>X"00",
30159=>X"00",
30160=>X"00",
30161=>X"00",
30162=>X"00",
30163=>X"00",
30164=>X"00",
30165=>X"00",
30166=>X"00",
30167=>X"00",
30168=>X"00",
30169=>X"00",
30170=>X"00",
30171=>X"00",
30172=>X"00",
30173=>X"00",
30174=>X"00",
30175=>X"00",
30176=>X"00",
30177=>X"00",
30178=>X"00",
30179=>X"00",
30180=>X"00",
30181=>X"00",
30182=>X"00",
30183=>X"00",
30184=>X"00",
30185=>X"00",
30186=>X"00",
30187=>X"00",
30188=>X"00",
30189=>X"00",
30190=>X"00",
30191=>X"00",
30192=>X"00",
30193=>X"00",
30194=>X"00",
30195=>X"00",
30196=>X"00",
30197=>X"00",
30198=>X"00",
30199=>X"00",
30200=>X"00",
30201=>X"00",
30202=>X"00",
30203=>X"00",
30204=>X"00",
30205=>X"00",
30206=>X"00",
30207=>X"00",
30208=>X"00",
30209=>X"00",
30210=>X"00",
30211=>X"00",
30212=>X"00",
30213=>X"00",
30214=>X"00",
30215=>X"00",
30216=>X"00",
30217=>X"00",
30218=>X"00",
30219=>X"00",
30220=>X"00",
30221=>X"00",
30222=>X"00",
30223=>X"00",
30224=>X"00",
30225=>X"00",
30226=>X"00",
30227=>X"00",
30228=>X"00",
30229=>X"00",
30230=>X"00",
30231=>X"00",
30232=>X"00",
30233=>X"00",
30234=>X"00",
30235=>X"00",
30236=>X"00",
30237=>X"00",
30238=>X"00",
30239=>X"00",
30240=>X"00",
30241=>X"00",
30242=>X"00",
30243=>X"00",
30244=>X"00",
30245=>X"00",
30246=>X"00",
30247=>X"00",
30248=>X"00",
30249=>X"00",
30250=>X"00",
30251=>X"00",
30252=>X"00",
30253=>X"00",
30254=>X"00",
30255=>X"00",
30256=>X"00",
30257=>X"00",
30258=>X"00",
30259=>X"00",
30260=>X"00",
30261=>X"00",
30262=>X"00",
30263=>X"00",
30264=>X"00",
30265=>X"00",
30266=>X"00",
30267=>X"00",
30268=>X"00",
30269=>X"00",
30270=>X"00",
30271=>X"00",
30272=>X"00",
30273=>X"00",
30274=>X"00",
30275=>X"00",
30276=>X"00",
30277=>X"00",
30278=>X"00",
30279=>X"00",
30280=>X"00",
30281=>X"00",
30282=>X"00",
30283=>X"00",
30284=>X"00",
30285=>X"00",
30286=>X"00",
30287=>X"00",
30288=>X"00",
30289=>X"00",
30290=>X"00",
30291=>X"00",
30292=>X"00",
30293=>X"00",
30294=>X"00",
30295=>X"00",
30296=>X"00",
30297=>X"00",
30298=>X"00",
30299=>X"00",
30300=>X"00",
30301=>X"00",
30302=>X"00",
30303=>X"00",
30304=>X"00",
30305=>X"00",
30306=>X"00",
30307=>X"00",
30308=>X"00",
30309=>X"00",
30310=>X"00",
30311=>X"00",
30312=>X"00",
30313=>X"00",
30314=>X"00",
30315=>X"00",
30316=>X"00",
30317=>X"00",
30318=>X"00",
30319=>X"00",
30320=>X"00",
30321=>X"00",
30322=>X"00",
30323=>X"00",
30324=>X"00",
30325=>X"00",
30326=>X"00",
30327=>X"00",
30328=>X"00",
30329=>X"00",
30330=>X"00",
30331=>X"00",
30332=>X"00",
30333=>X"00",
30334=>X"00",
30335=>X"00",
30336=>X"00",
30337=>X"00",
30338=>X"00",
30339=>X"00",
30340=>X"00",
30341=>X"00",
30342=>X"00",
30343=>X"00",
30344=>X"00",
30345=>X"00",
30346=>X"00",
30347=>X"00",
30348=>X"00",
30349=>X"00",
30350=>X"00",
30351=>X"00",
30352=>X"00",
30353=>X"00",
30354=>X"00",
30355=>X"00",
30356=>X"00",
30357=>X"00",
30358=>X"00",
30359=>X"00",
30360=>X"00",
30361=>X"00",
30362=>X"00",
30363=>X"00",
30364=>X"00",
30365=>X"00",
30366=>X"00",
30367=>X"00",
30368=>X"00",
30369=>X"00",
30370=>X"00",
30371=>X"00",
30372=>X"00",
30373=>X"00",
30374=>X"00",
30375=>X"00",
30376=>X"00",
30377=>X"00",
30378=>X"00",
30379=>X"00",
30380=>X"00",
30381=>X"00",
30382=>X"00",
30383=>X"00",
30384=>X"00",
30385=>X"00",
30386=>X"00",
30387=>X"00",
30388=>X"00",
30389=>X"00",
30390=>X"00",
30391=>X"00",
30392=>X"00",
30393=>X"00",
30394=>X"00",
30395=>X"00",
30396=>X"00",
30397=>X"00",
30398=>X"00",
30399=>X"00",
30400=>X"00",
30401=>X"00",
30402=>X"00",
30403=>X"00",
30404=>X"00",
30405=>X"00",
30406=>X"00",
30407=>X"00",
30408=>X"00",
30409=>X"00",
30410=>X"00",
30411=>X"00",
30412=>X"00",
30413=>X"00",
30414=>X"00",
30415=>X"00",
30416=>X"00",
30417=>X"00",
30418=>X"00",
30419=>X"00",
30420=>X"00",
30421=>X"00",
30422=>X"00",
30423=>X"00",
30424=>X"00",
30425=>X"00",
30426=>X"00",
30427=>X"00",
30428=>X"00",
30429=>X"00",
30430=>X"00",
30431=>X"00",
30432=>X"00",
30433=>X"00",
30434=>X"00",
30435=>X"00",
30436=>X"00",
30437=>X"00",
30438=>X"00",
30439=>X"00",
30440=>X"00",
30441=>X"00",
30442=>X"00",
30443=>X"00",
30444=>X"00",
30445=>X"00",
30446=>X"00",
30447=>X"00",
30448=>X"00",
30449=>X"00",
30450=>X"00",
30451=>X"00",
30452=>X"00",
30453=>X"00",
30454=>X"00",
30455=>X"00",
30456=>X"00",
30457=>X"00",
30458=>X"00",
30459=>X"00",
30460=>X"00",
30461=>X"00",
30462=>X"00",
30463=>X"00",
30464=>X"00",
30465=>X"00",
30466=>X"00",
30467=>X"00",
30468=>X"00",
30469=>X"00",
30470=>X"00",
30471=>X"00",
30472=>X"00",
30473=>X"00",
30474=>X"00",
30475=>X"00",
30476=>X"00",
30477=>X"00",
30478=>X"00",
30479=>X"00",
30480=>X"00",
30481=>X"00",
30482=>X"00",
30483=>X"00",
30484=>X"00",
30485=>X"00",
30486=>X"00",
30487=>X"00",
30488=>X"00",
30489=>X"00",
30490=>X"00",
30491=>X"00",
30492=>X"00",
30493=>X"00",
30494=>X"00",
30495=>X"00",
30496=>X"00",
30497=>X"00",
30498=>X"00",
30499=>X"00",
30500=>X"00",
30501=>X"00",
30502=>X"00",
30503=>X"00",
30504=>X"00",
30505=>X"00",
30506=>X"00",
30507=>X"00",
30508=>X"00",
30509=>X"00",
30510=>X"00",
30511=>X"00",
30512=>X"00",
30513=>X"00",
30514=>X"00",
30515=>X"00",
30516=>X"00",
30517=>X"00",
30518=>X"00",
30519=>X"00",
30520=>X"00",
30521=>X"00",
30522=>X"00",
30523=>X"00",
30524=>X"00",
30525=>X"00",
30526=>X"00",
30527=>X"00",
30528=>X"00",
30529=>X"00",
30530=>X"00",
30531=>X"00",
30532=>X"00",
30533=>X"00",
30534=>X"00",
30535=>X"00",
30536=>X"00",
30537=>X"00",
30538=>X"00",
30539=>X"00",
30540=>X"00",
30541=>X"00",
30542=>X"00",
30543=>X"00",
30544=>X"00",
30545=>X"00",
30546=>X"00",
30547=>X"00",
30548=>X"00",
30549=>X"00",
30550=>X"00",
30551=>X"00",
30552=>X"00",
30553=>X"00",
30554=>X"00",
30555=>X"00",
30556=>X"00",
30557=>X"00",
30558=>X"00",
30559=>X"00",
30560=>X"00",
30561=>X"00",
30562=>X"00",
30563=>X"00",
30564=>X"00",
30565=>X"00",
30566=>X"00",
30567=>X"00",
30568=>X"00",
30569=>X"00",
30570=>X"00",
30571=>X"00",
30572=>X"00",
30573=>X"00",
30574=>X"00",
30575=>X"00",
30576=>X"00",
30577=>X"00",
30578=>X"00",
30579=>X"00",
30580=>X"00",
30581=>X"00",
30582=>X"00",
30583=>X"00",
30584=>X"00",
30585=>X"00",
30586=>X"00",
30587=>X"00",
30588=>X"00",
30589=>X"00",
30590=>X"00",
30591=>X"00",
30592=>X"00",
30593=>X"00",
30594=>X"00",
30595=>X"00",
30596=>X"00",
30597=>X"00",
30598=>X"00",
30599=>X"00",
30600=>X"00",
30601=>X"00",
30602=>X"00",
30603=>X"00",
30604=>X"00",
30605=>X"00",
30606=>X"00",
30607=>X"00",
30608=>X"00",
30609=>X"00",
30610=>X"00",
30611=>X"00",
30612=>X"00",
30613=>X"00",
30614=>X"00",
30615=>X"00",
30616=>X"00",
30617=>X"00",
30618=>X"00",
30619=>X"00",
30620=>X"00",
30621=>X"00",
30622=>X"00",
30623=>X"00",
30624=>X"00",
30625=>X"00",
30626=>X"00",
30627=>X"00",
30628=>X"00",
30629=>X"00",
30630=>X"00",
30631=>X"00",
30632=>X"00",
30633=>X"00",
30634=>X"00",
30635=>X"00",
30636=>X"00",
30637=>X"00",
30638=>X"00",
30639=>X"00",
30640=>X"00",
30641=>X"00",
30642=>X"00",
30643=>X"00",
30644=>X"00",
30645=>X"00",
30646=>X"00",
30647=>X"00",
30648=>X"00",
30649=>X"00",
30650=>X"00",
30651=>X"00",
30652=>X"00",
30653=>X"00",
30654=>X"00",
30655=>X"00",
30656=>X"00",
30657=>X"00",
30658=>X"00",
30659=>X"00",
30660=>X"00",
30661=>X"00",
30662=>X"00",
30663=>X"00",
30664=>X"00",
30665=>X"00",
30666=>X"00",
30667=>X"00",
30668=>X"00",
30669=>X"00",
30670=>X"00",
30671=>X"00",
30672=>X"00",
30673=>X"00",
30674=>X"00",
30675=>X"00",
30676=>X"00",
30677=>X"00",
30678=>X"00",
30679=>X"00",
30680=>X"00",
30681=>X"00",
30682=>X"00",
30683=>X"00",
30684=>X"00",
30685=>X"00",
30686=>X"00",
30687=>X"00",
30688=>X"00",
30689=>X"00",
30690=>X"00",
30691=>X"00",
30692=>X"00",
30693=>X"00",
30694=>X"00",
30695=>X"00",
30696=>X"00",
30697=>X"00",
30698=>X"00",
30699=>X"00",
30700=>X"00",
30701=>X"00",
30702=>X"00",
30703=>X"00",
30704=>X"00",
30705=>X"00",
30706=>X"00",
30707=>X"00",
30708=>X"00",
30709=>X"00",
30710=>X"00",
30711=>X"00",
30712=>X"00",
30713=>X"00",
30714=>X"00",
30715=>X"00",
30716=>X"00",
30717=>X"00",
30718=>X"00",
30719=>X"00",
30720=>X"00",
30721=>X"00",
30722=>X"00",
30723=>X"00",
30724=>X"00",
30725=>X"00",
30726=>X"00",
30727=>X"00",
30728=>X"00",
30729=>X"00",
30730=>X"00",
30731=>X"00",
30732=>X"00",
30733=>X"00",
30734=>X"00",
30735=>X"00",
30736=>X"00",
30737=>X"00",
30738=>X"00",
30739=>X"00",
30740=>X"00",
30741=>X"00",
30742=>X"00",
30743=>X"00",
30744=>X"00",
30745=>X"00",
30746=>X"00",
30747=>X"00",
30748=>X"00",
30749=>X"00",
30750=>X"00",
30751=>X"00",
30752=>X"00",
30753=>X"00",
30754=>X"00",
30755=>X"00",
30756=>X"00",
30757=>X"00",
30758=>X"00",
30759=>X"00",
30760=>X"00",
30761=>X"00",
30762=>X"00",
30763=>X"00",
30764=>X"00",
30765=>X"00",
30766=>X"00",
30767=>X"00",
30768=>X"00",
30769=>X"00",
30770=>X"00",
30771=>X"00",
30772=>X"00",
30773=>X"00",
30774=>X"00",
30775=>X"00",
30776=>X"00",
30777=>X"00",
30778=>X"00",
30779=>X"00",
30780=>X"00",
30781=>X"00",
30782=>X"00",
30783=>X"00",
30784=>X"00",
30785=>X"00",
30786=>X"00",
30787=>X"00",
30788=>X"00",
30789=>X"00",
30790=>X"00",
30791=>X"00",
30792=>X"00",
30793=>X"00",
30794=>X"00",
30795=>X"00",
30796=>X"00",
30797=>X"00",
30798=>X"00",
30799=>X"00",
30800=>X"00",
30801=>X"00",
30802=>X"00",
30803=>X"00",
30804=>X"00",
30805=>X"00",
30806=>X"00",
30807=>X"00",
30808=>X"00",
30809=>X"00",
30810=>X"00",
30811=>X"00",
30812=>X"00",
30813=>X"00",
30814=>X"00",
30815=>X"00",
30816=>X"00",
30817=>X"00",
30818=>X"00",
30819=>X"00",
30820=>X"00",
30821=>X"00",
30822=>X"00",
30823=>X"00",
30824=>X"00",
30825=>X"00",
30826=>X"00",
30827=>X"00",
30828=>X"00",
30829=>X"00",
30830=>X"00",
30831=>X"00",
30832=>X"00",
30833=>X"00",
30834=>X"00",
30835=>X"00",
30836=>X"00",
30837=>X"00",
30838=>X"00",
30839=>X"00",
30840=>X"00",
30841=>X"00",
30842=>X"00",
30843=>X"00",
30844=>X"00",
30845=>X"00",
30846=>X"00",
30847=>X"00",
30848=>X"00",
30849=>X"00",
30850=>X"00",
30851=>X"00",
30852=>X"00",
30853=>X"00",
30854=>X"00",
30855=>X"00",
30856=>X"00",
30857=>X"00",
30858=>X"00",
30859=>X"00",
30860=>X"00",
30861=>X"00",
30862=>X"00",
30863=>X"00",
30864=>X"00",
30865=>X"00",
30866=>X"00",
30867=>X"00",
30868=>X"00",
30869=>X"00",
30870=>X"00",
30871=>X"00",
30872=>X"00",
30873=>X"00",
30874=>X"00",
30875=>X"00",
30876=>X"00",
30877=>X"00",
30878=>X"00",
30879=>X"00",
30880=>X"00",
30881=>X"00",
30882=>X"00",
30883=>X"00",
30884=>X"00",
30885=>X"00",
30886=>X"00",
30887=>X"00",
30888=>X"00",
30889=>X"00",
30890=>X"00",
30891=>X"00",
30892=>X"00",
30893=>X"00",
30894=>X"00",
30895=>X"00",
30896=>X"00",
30897=>X"00",
30898=>X"00",
30899=>X"00",
30900=>X"00",
30901=>X"00",
30902=>X"00",
30903=>X"00",
30904=>X"00",
30905=>X"00",
30906=>X"00",
30907=>X"00",
30908=>X"00",
30909=>X"00",
30910=>X"00",
30911=>X"00",
30912=>X"00",
30913=>X"00",
30914=>X"00",
30915=>X"00",
30916=>X"00",
30917=>X"00",
30918=>X"00",
30919=>X"00",
30920=>X"00",
30921=>X"00",
30922=>X"00",
30923=>X"00",
30924=>X"00",
30925=>X"00",
30926=>X"00",
30927=>X"00",
30928=>X"00",
30929=>X"00",
30930=>X"00",
30931=>X"00",
30932=>X"00",
30933=>X"00",
30934=>X"00",
30935=>X"00",
30936=>X"00",
30937=>X"00",
30938=>X"00",
30939=>X"00",
30940=>X"00",
30941=>X"00",
30942=>X"00",
30943=>X"00",
30944=>X"00",
30945=>X"00",
30946=>X"00",
30947=>X"00",
30948=>X"00",
30949=>X"00",
30950=>X"00",
30951=>X"00",
30952=>X"00",
30953=>X"00",
30954=>X"00",
30955=>X"00",
30956=>X"00",
30957=>X"00",
30958=>X"00",
30959=>X"00",
30960=>X"00",
30961=>X"00",
30962=>X"00",
30963=>X"00",
30964=>X"00",
30965=>X"00",
30966=>X"00",
30967=>X"00",
30968=>X"00",
30969=>X"00",
30970=>X"00",
30971=>X"00",
30972=>X"00",
30973=>X"00",
30974=>X"00",
30975=>X"00",
30976=>X"00",
30977=>X"00",
30978=>X"00",
30979=>X"00",
30980=>X"00",
30981=>X"00",
30982=>X"00",
30983=>X"00",
30984=>X"00",
30985=>X"00",
30986=>X"00",
30987=>X"00",
30988=>X"00",
30989=>X"00",
30990=>X"00",
30991=>X"00",
30992=>X"00",
30993=>X"00",
30994=>X"00",
30995=>X"00",
30996=>X"00",
30997=>X"00",
30998=>X"00",
30999=>X"00",
31000=>X"00",
31001=>X"00",
31002=>X"00",
31003=>X"00",
31004=>X"00",
31005=>X"00",
31006=>X"00",
31007=>X"00",
31008=>X"00",
31009=>X"00",
31010=>X"00",
31011=>X"00",
31012=>X"00",
31013=>X"00",
31014=>X"00",
31015=>X"00",
31016=>X"00",
31017=>X"00",
31018=>X"00",
31019=>X"00",
31020=>X"00",
31021=>X"00",
31022=>X"00",
31023=>X"00",
31024=>X"00",
31025=>X"00",
31026=>X"00",
31027=>X"00",
31028=>X"00",
31029=>X"00",
31030=>X"00",
31031=>X"00",
31032=>X"00",
31033=>X"00",
31034=>X"00",
31035=>X"00",
31036=>X"00",
31037=>X"00",
31038=>X"00",
31039=>X"00",
31040=>X"00",
31041=>X"00",
31042=>X"00",
31043=>X"00",
31044=>X"00",
31045=>X"00",
31046=>X"00",
31047=>X"00",
31048=>X"00",
31049=>X"00",
31050=>X"00",
31051=>X"00",
31052=>X"00",
31053=>X"00",
31054=>X"00",
31055=>X"00",
31056=>X"00",
31057=>X"00",
31058=>X"00",
31059=>X"00",
31060=>X"00",
31061=>X"00",
31062=>X"00",
31063=>X"00",
31064=>X"00",
31065=>X"00",
31066=>X"00",
31067=>X"00",
31068=>X"00",
31069=>X"00",
31070=>X"00",
31071=>X"00",
31072=>X"00",
31073=>X"00",
31074=>X"00",
31075=>X"00",
31076=>X"00",
31077=>X"00",
31078=>X"00",
31079=>X"00",
31080=>X"00",
31081=>X"00",
31082=>X"00",
31083=>X"00",
31084=>X"00",
31085=>X"00",
31086=>X"00",
31087=>X"00",
31088=>X"00",
31089=>X"00",
31090=>X"00",
31091=>X"00",
31092=>X"00",
31093=>X"00",
31094=>X"00",
31095=>X"00",
31096=>X"00",
31097=>X"00",
31098=>X"00",
31099=>X"00",
31100=>X"00",
31101=>X"00",
31102=>X"00",
31103=>X"00",
31104=>X"00",
31105=>X"00",
31106=>X"00",
31107=>X"00",
31108=>X"00",
31109=>X"00",
31110=>X"00",
31111=>X"00",
31112=>X"00",
31113=>X"00",
31114=>X"00",
31115=>X"00",
31116=>X"00",
31117=>X"00",
31118=>X"00",
31119=>X"00",
31120=>X"00",
31121=>X"00",
31122=>X"00",
31123=>X"00",
31124=>X"00",
31125=>X"00",
31126=>X"00",
31127=>X"00",
31128=>X"00",
31129=>X"00",
31130=>X"00",
31131=>X"00",
31132=>X"00",
31133=>X"00",
31134=>X"00",
31135=>X"00",
31136=>X"00",
31137=>X"00",
31138=>X"00",
31139=>X"00",
31140=>X"00",
31141=>X"00",
31142=>X"00",
31143=>X"00",
31144=>X"00",
31145=>X"00",
31146=>X"00",
31147=>X"00",
31148=>X"00",
31149=>X"00",
31150=>X"00",
31151=>X"00",
31152=>X"00",
31153=>X"00",
31154=>X"00",
31155=>X"00",
31156=>X"00",
31157=>X"00",
31158=>X"00",
31159=>X"00",
31160=>X"00",
31161=>X"00",
31162=>X"00",
31163=>X"00",
31164=>X"00",
31165=>X"00",
31166=>X"00",
31167=>X"00",
31168=>X"00",
31169=>X"00",
31170=>X"00",
31171=>X"00",
31172=>X"00",
31173=>X"00",
31174=>X"00",
31175=>X"00",
31176=>X"00",
31177=>X"00",
31178=>X"00",
31179=>X"00",
31180=>X"00",
31181=>X"00",
31182=>X"00",
31183=>X"00",
31184=>X"00",
31185=>X"00",
31186=>X"00",
31187=>X"00",
31188=>X"00",
31189=>X"00",
31190=>X"00",
31191=>X"00",
31192=>X"00",
31193=>X"00",
31194=>X"00",
31195=>X"00",
31196=>X"00",
31197=>X"00",
31198=>X"00",
31199=>X"00",
31200=>X"00",
31201=>X"00",
31202=>X"00",
31203=>X"00",
31204=>X"00",
31205=>X"00",
31206=>X"00",
31207=>X"00",
31208=>X"00",
31209=>X"00",
31210=>X"00",
31211=>X"00",
31212=>X"00",
31213=>X"00",
31214=>X"00",
31215=>X"00",
31216=>X"00",
31217=>X"00",
31218=>X"00",
31219=>X"00",
31220=>X"00",
31221=>X"00",
31222=>X"00",
31223=>X"00",
31224=>X"00",
31225=>X"00",
31226=>X"00",
31227=>X"00",
31228=>X"00",
31229=>X"00",
31230=>X"00",
31231=>X"00",
31232=>X"00",
31233=>X"00",
31234=>X"00",
31235=>X"00",
31236=>X"00",
31237=>X"00",
31238=>X"00",
31239=>X"00",
31240=>X"00",
31241=>X"00",
31242=>X"00",
31243=>X"00",
31244=>X"00",
31245=>X"00",
31246=>X"00",
31247=>X"00",
31248=>X"00",
31249=>X"00",
31250=>X"00",
31251=>X"00",
31252=>X"00",
31253=>X"00",
31254=>X"00",
31255=>X"00",
31256=>X"00",
31257=>X"00",
31258=>X"00",
31259=>X"00",
31260=>X"00",
31261=>X"00",
31262=>X"00",
31263=>X"00",
31264=>X"00",
31265=>X"00",
31266=>X"00",
31267=>X"00",
31268=>X"00",
31269=>X"00",
31270=>X"00",
31271=>X"00",
31272=>X"00",
31273=>X"00",
31274=>X"00",
31275=>X"00",
31276=>X"00",
31277=>X"00",
31278=>X"00",
31279=>X"00",
31280=>X"00",
31281=>X"00",
31282=>X"00",
31283=>X"00",
31284=>X"00",
31285=>X"00",
31286=>X"00",
31287=>X"00",
31288=>X"00",
31289=>X"00",
31290=>X"00",
31291=>X"00",
31292=>X"00",
31293=>X"00",
31294=>X"00",
31295=>X"00",
31296=>X"00",
31297=>X"00",
31298=>X"00",
31299=>X"00",
31300=>X"00",
31301=>X"00",
31302=>X"00",
31303=>X"00",
31304=>X"00",
31305=>X"00",
31306=>X"00",
31307=>X"00",
31308=>X"00",
31309=>X"00",
31310=>X"00",
31311=>X"00",
31312=>X"00",
31313=>X"00",
31314=>X"00",
31315=>X"00",
31316=>X"00",
31317=>X"00",
31318=>X"00",
31319=>X"00",
31320=>X"00",
31321=>X"00",
31322=>X"00",
31323=>X"00",
31324=>X"00",
31325=>X"00",
31326=>X"00",
31327=>X"00",
31328=>X"00",
31329=>X"00",
31330=>X"00",
31331=>X"00",
31332=>X"00",
31333=>X"00",
31334=>X"00",
31335=>X"00",
31336=>X"00",
31337=>X"00",
31338=>X"00",
31339=>X"00",
31340=>X"00",
31341=>X"00",
31342=>X"00",
31343=>X"00",
31344=>X"00",
31345=>X"00",
31346=>X"00",
31347=>X"00",
31348=>X"00",
31349=>X"00",
31350=>X"00",
31351=>X"00",
31352=>X"00",
31353=>X"00",
31354=>X"00",
31355=>X"00",
31356=>X"00",
31357=>X"00",
31358=>X"00",
31359=>X"00",
31360=>X"00",
31361=>X"00",
31362=>X"00",
31363=>X"00",
31364=>X"00",
31365=>X"00",
31366=>X"00",
31367=>X"00",
31368=>X"00",
31369=>X"00",
31370=>X"00",
31371=>X"00",
31372=>X"00",
31373=>X"00",
31374=>X"00",
31375=>X"00",
31376=>X"00",
31377=>X"00",
31378=>X"00",
31379=>X"00",
31380=>X"00",
31381=>X"00",
31382=>X"00",
31383=>X"00",
31384=>X"00",
31385=>X"00",
31386=>X"00",
31387=>X"00",
31388=>X"00",
31389=>X"00",
31390=>X"00",
31391=>X"00",
31392=>X"00",
31393=>X"00",
31394=>X"00",
31395=>X"00",
31396=>X"00",
31397=>X"00",
31398=>X"00",
31399=>X"00",
31400=>X"00",
31401=>X"00",
31402=>X"00",
31403=>X"00",
31404=>X"00",
31405=>X"00",
31406=>X"00",
31407=>X"00",
31408=>X"00",
31409=>X"00",
31410=>X"00",
31411=>X"00",
31412=>X"00",
31413=>X"00",
31414=>X"00",
31415=>X"00",
31416=>X"00",
31417=>X"00",
31418=>X"00",
31419=>X"00",
31420=>X"00",
31421=>X"00",
31422=>X"00",
31423=>X"00",
31424=>X"00",
31425=>X"00",
31426=>X"00",
31427=>X"00",
31428=>X"00",
31429=>X"00",
31430=>X"00",
31431=>X"00",
31432=>X"00",
31433=>X"00",
31434=>X"00",
31435=>X"00",
31436=>X"00",
31437=>X"00",
31438=>X"00",
31439=>X"00",
31440=>X"00",
31441=>X"00",
31442=>X"00",
31443=>X"00",
31444=>X"00",
31445=>X"00",
31446=>X"00",
31447=>X"00",
31448=>X"00",
31449=>X"00",
31450=>X"00",
31451=>X"00",
31452=>X"00",
31453=>X"00",
31454=>X"00",
31455=>X"00",
31456=>X"00",
31457=>X"00",
31458=>X"00",
31459=>X"00",
31460=>X"00",
31461=>X"00",
31462=>X"00",
31463=>X"00",
31464=>X"00",
31465=>X"00",
31466=>X"00",
31467=>X"00",
31468=>X"00",
31469=>X"00",
31470=>X"00",
31471=>X"00",
31472=>X"00",
31473=>X"00",
31474=>X"00",
31475=>X"00",
31476=>X"00",
31477=>X"00",
31478=>X"00",
31479=>X"00",
31480=>X"00",
31481=>X"00",
31482=>X"00",
31483=>X"00",
31484=>X"00",
31485=>X"00",
31486=>X"00",
31487=>X"00",
31488=>X"00",
31489=>X"00",
31490=>X"00",
31491=>X"00",
31492=>X"00",
31493=>X"00",
31494=>X"00",
31495=>X"00",
31496=>X"00",
31497=>X"00",
31498=>X"00",
31499=>X"00",
31500=>X"00",
31501=>X"00",
31502=>X"00",
31503=>X"00",
31504=>X"00",
31505=>X"00",
31506=>X"00",
31507=>X"00",
31508=>X"00",
31509=>X"00",
31510=>X"00",
31511=>X"00",
31512=>X"00",
31513=>X"00",
31514=>X"00",
31515=>X"00",
31516=>X"00",
31517=>X"00",
31518=>X"00",
31519=>X"00",
31520=>X"00",
31521=>X"00",
31522=>X"00",
31523=>X"00",
31524=>X"00",
31525=>X"00",
31526=>X"00",
31527=>X"00",
31528=>X"00",
31529=>X"00",
31530=>X"00",
31531=>X"00",
31532=>X"00",
31533=>X"00",
31534=>X"00",
31535=>X"00",
31536=>X"00",
31537=>X"00",
31538=>X"00",
31539=>X"00",
31540=>X"00",
31541=>X"00",
31542=>X"00",
31543=>X"00",
31544=>X"00",
31545=>X"00",
31546=>X"00",
31547=>X"00",
31548=>X"00",
31549=>X"00",
31550=>X"00",
31551=>X"00",
31552=>X"00",
31553=>X"00",
31554=>X"00",
31555=>X"00",
31556=>X"00",
31557=>X"00",
31558=>X"00",
31559=>X"00",
31560=>X"00",
31561=>X"00",
31562=>X"00",
31563=>X"00",
31564=>X"00",
31565=>X"00",
31566=>X"00",
31567=>X"00",
31568=>X"00",
31569=>X"00",
31570=>X"00",
31571=>X"00",
31572=>X"00",
31573=>X"00",
31574=>X"00",
31575=>X"00",
31576=>X"00",
31577=>X"00",
31578=>X"00",
31579=>X"00",
31580=>X"00",
31581=>X"00",
31582=>X"00",
31583=>X"00",
31584=>X"00",
31585=>X"00",
31586=>X"00",
31587=>X"00",
31588=>X"00",
31589=>X"00",
31590=>X"00",
31591=>X"00",
31592=>X"00",
31593=>X"00",
31594=>X"00",
31595=>X"00",
31596=>X"00",
31597=>X"00",
31598=>X"00",
31599=>X"00",
31600=>X"00",
31601=>X"00",
31602=>X"00",
31603=>X"00",
31604=>X"00",
31605=>X"00",
31606=>X"00",
31607=>X"00",
31608=>X"00",
31609=>X"00",
31610=>X"00",
31611=>X"00",
31612=>X"00",
31613=>X"00",
31614=>X"00",
31615=>X"00",
31616=>X"00",
31617=>X"00",
31618=>X"00",
31619=>X"00",
31620=>X"00",
31621=>X"00",
31622=>X"00",
31623=>X"00",
31624=>X"00",
31625=>X"00",
31626=>X"00",
31627=>X"00",
31628=>X"00",
31629=>X"00",
31630=>X"00",
31631=>X"00",
31632=>X"00",
31633=>X"00",
31634=>X"00",
31635=>X"00",
31636=>X"00",
31637=>X"00",
31638=>X"00",
31639=>X"00",
31640=>X"00",
31641=>X"00",
31642=>X"00",
31643=>X"00",
31644=>X"00",
31645=>X"00",
31646=>X"00",
31647=>X"00",
31648=>X"00",
31649=>X"00",
31650=>X"00",
31651=>X"00",
31652=>X"00",
31653=>X"00",
31654=>X"00",
31655=>X"00",
31656=>X"00",
31657=>X"00",
31658=>X"00",
31659=>X"00",
31660=>X"00",
31661=>X"00",
31662=>X"00",
31663=>X"00",
31664=>X"00",
31665=>X"00",
31666=>X"00",
31667=>X"00",
31668=>X"00",
31669=>X"00",
31670=>X"00",
31671=>X"00",
31672=>X"00",
31673=>X"00",
31674=>X"00",
31675=>X"00",
31676=>X"00",
31677=>X"00",
31678=>X"00",
31679=>X"00",
31680=>X"00",
31681=>X"00",
31682=>X"00",
31683=>X"00",
31684=>X"00",
31685=>X"00",
31686=>X"00",
31687=>X"00",
31688=>X"00",
31689=>X"00",
31690=>X"00",
31691=>X"00",
31692=>X"00",
31693=>X"00",
31694=>X"00",
31695=>X"00",
31696=>X"00",
31697=>X"00",
31698=>X"00",
31699=>X"00",
31700=>X"00",
31701=>X"00",
31702=>X"00",
31703=>X"00",
31704=>X"00",
31705=>X"00",
31706=>X"00",
31707=>X"00",
31708=>X"00",
31709=>X"00",
31710=>X"00",
31711=>X"00",
31712=>X"00",
31713=>X"00",
31714=>X"00",
31715=>X"00",
31716=>X"00",
31717=>X"00",
31718=>X"00",
31719=>X"00",
31720=>X"00",
31721=>X"00",
31722=>X"00",
31723=>X"00",
31724=>X"00",
31725=>X"00",
31726=>X"00",
31727=>X"00",
31728=>X"00",
31729=>X"00",
31730=>X"00",
31731=>X"00",
31732=>X"00",
31733=>X"00",
31734=>X"00",
31735=>X"00",
31736=>X"00",
31737=>X"00",
31738=>X"00",
31739=>X"00",
31740=>X"00",
31741=>X"00",
31742=>X"00",
31743=>X"00",
31744=>X"00",
31745=>X"00",
31746=>X"00",
31747=>X"00",
31748=>X"00",
31749=>X"00",
31750=>X"00",
31751=>X"00",
31752=>X"00",
31753=>X"00",
31754=>X"00",
31755=>X"00",
31756=>X"00",
31757=>X"00",
31758=>X"00",
31759=>X"00",
31760=>X"00",
31761=>X"00",
31762=>X"00",
31763=>X"00",
31764=>X"00",
31765=>X"00",
31766=>X"00",
31767=>X"00",
31768=>X"00",
31769=>X"00",
31770=>X"00",
31771=>X"00",
31772=>X"00",
31773=>X"00",
31774=>X"00",
31775=>X"00",
31776=>X"00",
31777=>X"00",
31778=>X"00",
31779=>X"00",
31780=>X"00",
31781=>X"00",
31782=>X"00",
31783=>X"00",
31784=>X"00",
31785=>X"00",
31786=>X"00",
31787=>X"00",
31788=>X"00",
31789=>X"00",
31790=>X"00",
31791=>X"00",
31792=>X"00",
31793=>X"00",
31794=>X"00",
31795=>X"00",
31796=>X"00",
31797=>X"00",
31798=>X"00",
31799=>X"00",
31800=>X"00",
31801=>X"00",
31802=>X"00",
31803=>X"00",
31804=>X"00",
31805=>X"00",
31806=>X"00",
31807=>X"00",
31808=>X"00",
31809=>X"00",
31810=>X"00",
31811=>X"00",
31812=>X"00",
31813=>X"00",
31814=>X"00",
31815=>X"00",
31816=>X"00",
31817=>X"00",
31818=>X"00",
31819=>X"00",
31820=>X"00",
31821=>X"00",
31822=>X"00",
31823=>X"00",
31824=>X"00",
31825=>X"00",
31826=>X"00",
31827=>X"00",
31828=>X"00",
31829=>X"00",
31830=>X"00",
31831=>X"00",
31832=>X"00",
31833=>X"00",
31834=>X"00",
31835=>X"00",
31836=>X"00",
31837=>X"00",
31838=>X"00",
31839=>X"00",
31840=>X"00",
31841=>X"00",
31842=>X"00",
31843=>X"00",
31844=>X"00",
31845=>X"00",
31846=>X"00",
31847=>X"00",
31848=>X"00",
31849=>X"00",
31850=>X"00",
31851=>X"00",
31852=>X"00",
31853=>X"00",
31854=>X"00",
31855=>X"00",
31856=>X"00",
31857=>X"00",
31858=>X"00",
31859=>X"00",
31860=>X"00",
31861=>X"00",
31862=>X"00",
31863=>X"00",
31864=>X"00",
31865=>X"00",
31866=>X"00",
31867=>X"00",
31868=>X"00",
31869=>X"00",
31870=>X"00",
31871=>X"00",
31872=>X"00",
31873=>X"00",
31874=>X"00",
31875=>X"00",
31876=>X"00",
31877=>X"00",
31878=>X"00",
31879=>X"00",
31880=>X"00",
31881=>X"00",
31882=>X"00",
31883=>X"00",
31884=>X"00",
31885=>X"00",
31886=>X"00",
31887=>X"00",
31888=>X"00",
31889=>X"00",
31890=>X"00",
31891=>X"00",
31892=>X"00",
31893=>X"00",
31894=>X"00",
31895=>X"00",
31896=>X"00",
31897=>X"00",
31898=>X"00",
31899=>X"00",
31900=>X"00",
31901=>X"00",
31902=>X"00",
31903=>X"00",
31904=>X"00",
31905=>X"00",
31906=>X"00",
31907=>X"00",
31908=>X"00",
31909=>X"00",
31910=>X"00",
31911=>X"00",
31912=>X"00",
31913=>X"00",
31914=>X"00",
31915=>X"00",
31916=>X"00",
31917=>X"00",
31918=>X"00",
31919=>X"00",
31920=>X"00",
31921=>X"00",
31922=>X"00",
31923=>X"00",
31924=>X"00",
31925=>X"00",
31926=>X"00",
31927=>X"00",
31928=>X"00",
31929=>X"00",
31930=>X"00",
31931=>X"00",
31932=>X"00",
31933=>X"00",
31934=>X"00",
31935=>X"00",
31936=>X"00",
31937=>X"00",
31938=>X"00",
31939=>X"00",
31940=>X"00",
31941=>X"00",
31942=>X"00",
31943=>X"00",
31944=>X"00",
31945=>X"00",
31946=>X"00",
31947=>X"00",
31948=>X"00",
31949=>X"00",
31950=>X"00",
31951=>X"00",
31952=>X"00",
31953=>X"00",
31954=>X"00",
31955=>X"00",
31956=>X"00",
31957=>X"00",
31958=>X"00",
31959=>X"00",
31960=>X"00",
31961=>X"00",
31962=>X"00",
31963=>X"00",
31964=>X"00",
31965=>X"00",
31966=>X"00",
31967=>X"00",
31968=>X"00",
31969=>X"00",
31970=>X"00",
31971=>X"00",
31972=>X"00",
31973=>X"00",
31974=>X"00",
31975=>X"00",
31976=>X"00",
31977=>X"00",
31978=>X"00",
31979=>X"00",
31980=>X"00",
31981=>X"00",
31982=>X"00",
31983=>X"00",
31984=>X"00",
31985=>X"00",
31986=>X"00",
31987=>X"00",
31988=>X"00",
31989=>X"00",
31990=>X"00",
31991=>X"00",
31992=>X"00",
31993=>X"00",
31994=>X"00",
31995=>X"00",
31996=>X"00",
31997=>X"00",
31998=>X"00",
31999=>X"00",
32000=>X"00",
32001=>X"00",
32002=>X"00",
32003=>X"00",
32004=>X"00",
32005=>X"00",
32006=>X"00",
32007=>X"00",
32008=>X"00",
32009=>X"00",
32010=>X"00",
32011=>X"00",
32012=>X"00",
32013=>X"00",
32014=>X"00",
32015=>X"00",
32016=>X"00",
32017=>X"00",
32018=>X"00",
32019=>X"00",
32020=>X"00",
32021=>X"00",
32022=>X"00",
32023=>X"00",
32024=>X"00",
32025=>X"00",
32026=>X"00",
32027=>X"00",
32028=>X"00",
32029=>X"00",
32030=>X"00",
32031=>X"00",
32032=>X"00",
32033=>X"00",
32034=>X"00",
32035=>X"00",
32036=>X"00",
32037=>X"00",
32038=>X"00",
32039=>X"00",
32040=>X"00",
32041=>X"00",
32042=>X"00",
32043=>X"00",
32044=>X"00",
32045=>X"00",
32046=>X"00",
32047=>X"00",
32048=>X"00",
32049=>X"00",
32050=>X"00",
32051=>X"00",
32052=>X"00",
32053=>X"00",
32054=>X"00",
32055=>X"00",
32056=>X"00",
32057=>X"00",
32058=>X"00",
32059=>X"00",
32060=>X"00",
32061=>X"00",
32062=>X"00",
32063=>X"00",
32064=>X"00",
32065=>X"00",
32066=>X"00",
32067=>X"00",
32068=>X"00",
32069=>X"00",
32070=>X"00",
32071=>X"00",
32072=>X"00",
32073=>X"00",
32074=>X"00",
32075=>X"00",
32076=>X"00",
32077=>X"00",
32078=>X"00",
32079=>X"00",
32080=>X"00",
32081=>X"00",
32082=>X"00",
32083=>X"00",
32084=>X"00",
32085=>X"00",
32086=>X"00",
32087=>X"00",
32088=>X"00",
32089=>X"00",
32090=>X"00",
32091=>X"00",
32092=>X"00",
32093=>X"00",
32094=>X"00",
32095=>X"00",
32096=>X"00",
32097=>X"00",
32098=>X"00",
32099=>X"00",
32100=>X"00",
32101=>X"00",
32102=>X"00",
32103=>X"00",
32104=>X"00",
32105=>X"00",
32106=>X"00",
32107=>X"00",
32108=>X"00",
32109=>X"00",
32110=>X"00",
32111=>X"00",
32112=>X"00",
32113=>X"00",
32114=>X"00",
32115=>X"00",
32116=>X"00",
32117=>X"00",
32118=>X"00",
32119=>X"00",
32120=>X"00",
32121=>X"00",
32122=>X"00",
32123=>X"00",
32124=>X"00",
32125=>X"00",
32126=>X"00",
32127=>X"00",
32128=>X"00",
32129=>X"00",
32130=>X"00",
32131=>X"00",
32132=>X"00",
32133=>X"00",
32134=>X"00",
32135=>X"00",
32136=>X"00",
32137=>X"00",
32138=>X"00",
32139=>X"00",
32140=>X"00",
32141=>X"00",
32142=>X"00",
32143=>X"00",
32144=>X"00",
32145=>X"00",
32146=>X"00",
32147=>X"00",
32148=>X"00",
32149=>X"00",
32150=>X"00",
32151=>X"00",
32152=>X"00",
32153=>X"00",
32154=>X"00",
32155=>X"00",
32156=>X"00",
32157=>X"00",
32158=>X"00",
32159=>X"00",
32160=>X"00",
32161=>X"00",
32162=>X"00",
32163=>X"00",
32164=>X"00",
32165=>X"00",
32166=>X"00",
32167=>X"00",
32168=>X"00",
32169=>X"00",
32170=>X"00",
32171=>X"00",
32172=>X"00",
32173=>X"00",
32174=>X"00",
32175=>X"00",
32176=>X"00",
32177=>X"00",
32178=>X"00",
32179=>X"00",
32180=>X"00",
32181=>X"00",
32182=>X"00",
32183=>X"00",
32184=>X"00",
32185=>X"00",
32186=>X"00",
32187=>X"00",
32188=>X"00",
32189=>X"00",
32190=>X"00",
32191=>X"00",
32192=>X"00",
32193=>X"00",
32194=>X"00",
32195=>X"00",
32196=>X"00",
32197=>X"00",
32198=>X"00",
32199=>X"00",
32200=>X"00",
32201=>X"00",
32202=>X"00",
32203=>X"00",
32204=>X"00",
32205=>X"00",
32206=>X"00",
32207=>X"00",
32208=>X"00",
32209=>X"00",
32210=>X"00",
32211=>X"00",
32212=>X"00",
32213=>X"00",
32214=>X"00",
32215=>X"00",
32216=>X"00",
32217=>X"00",
32218=>X"00",
32219=>X"00",
32220=>X"00",
32221=>X"00",
32222=>X"00",
32223=>X"00",
32224=>X"00",
32225=>X"00",
32226=>X"00",
32227=>X"00",
32228=>X"00",
32229=>X"00",
32230=>X"00",
32231=>X"00",
32232=>X"00",
32233=>X"00",
32234=>X"00",
32235=>X"00",
32236=>X"00",
32237=>X"00",
32238=>X"00",
32239=>X"00",
32240=>X"00",
32241=>X"00",
32242=>X"00",
32243=>X"00",
32244=>X"00",
32245=>X"00",
32246=>X"00",
32247=>X"00",
32248=>X"00",
32249=>X"00",
32250=>X"00",
32251=>X"00",
32252=>X"00",
32253=>X"00",
32254=>X"00",
32255=>X"00",
32256=>X"00",
32257=>X"00",
32258=>X"00",
32259=>X"00",
32260=>X"00",
32261=>X"00",
32262=>X"00",
32263=>X"00",
32264=>X"00",
32265=>X"00",
32266=>X"00",
32267=>X"00",
32268=>X"00",
32269=>X"00",
32270=>X"00",
32271=>X"00",
32272=>X"00",
32273=>X"00",
32274=>X"00",
32275=>X"00",
32276=>X"00",
32277=>X"00",
32278=>X"00",
32279=>X"00",
32280=>X"00",
32281=>X"00",
32282=>X"00",
32283=>X"00",
32284=>X"00",
32285=>X"00",
32286=>X"00",
32287=>X"00",
32288=>X"00",
32289=>X"00",
32290=>X"00",
32291=>X"00",
32292=>X"00",
32293=>X"00",
32294=>X"00",
32295=>X"00",
32296=>X"00",
32297=>X"00",
32298=>X"00",
32299=>X"00",
32300=>X"00",
32301=>X"00",
32302=>X"00",
32303=>X"00",
32304=>X"00",
32305=>X"00",
32306=>X"00",
32307=>X"00",
32308=>X"00",
32309=>X"00",
32310=>X"00",
32311=>X"00",
32312=>X"00",
32313=>X"00",
32314=>X"00",
32315=>X"00",
32316=>X"00",
32317=>X"00",
32318=>X"00",
32319=>X"00",
32320=>X"00",
32321=>X"00",
32322=>X"00",
32323=>X"00",
32324=>X"00",
32325=>X"00",
32326=>X"00",
32327=>X"00",
32328=>X"00",
32329=>X"00",
32330=>X"00",
32331=>X"00",
32332=>X"00",
32333=>X"00",
32334=>X"00",
32335=>X"00",
32336=>X"00",
32337=>X"00",
32338=>X"00",
32339=>X"00",
32340=>X"00",
32341=>X"00",
32342=>X"00",
32343=>X"00",
32344=>X"00",
32345=>X"00",
32346=>X"00",
32347=>X"00",
32348=>X"00",
32349=>X"00",
32350=>X"00",
32351=>X"00",
32352=>X"00",
32353=>X"00",
32354=>X"00",
32355=>X"00",
32356=>X"00",
32357=>X"00",
32358=>X"00",
32359=>X"00",
32360=>X"00",
32361=>X"00",
32362=>X"00",
32363=>X"00",
32364=>X"00",
32365=>X"00",
32366=>X"00",
32367=>X"00",
32368=>X"00",
32369=>X"00",
32370=>X"00",
32371=>X"00",
32372=>X"00",
32373=>X"00",
32374=>X"00",
32375=>X"00",
32376=>X"00",
32377=>X"00",
32378=>X"00",
32379=>X"00",
32380=>X"00",
32381=>X"00",
32382=>X"00",
32383=>X"00",
32384=>X"00",
32385=>X"00",
32386=>X"00",
32387=>X"00",
32388=>X"00",
32389=>X"00",
32390=>X"00",
32391=>X"00",
32392=>X"00",
32393=>X"00",
32394=>X"00",
32395=>X"00",
32396=>X"00",
32397=>X"00",
32398=>X"00",
32399=>X"00",
32400=>X"00",
32401=>X"00",
32402=>X"00",
32403=>X"00",
32404=>X"00",
32405=>X"00",
32406=>X"00",
32407=>X"00",
32408=>X"00",
32409=>X"00",
32410=>X"00",
32411=>X"00",
32412=>X"00",
32413=>X"00",
32414=>X"00",
32415=>X"00",
32416=>X"00",
32417=>X"00",
32418=>X"00",
32419=>X"00",
32420=>X"00",
32421=>X"00",
32422=>X"00",
32423=>X"00",
32424=>X"00",
32425=>X"00",
32426=>X"00",
32427=>X"00",
32428=>X"00",
32429=>X"00",
32430=>X"00",
32431=>X"00",
32432=>X"00",
32433=>X"00",
32434=>X"00",
32435=>X"00",
32436=>X"00",
32437=>X"00",
32438=>X"00",
32439=>X"00",
32440=>X"00",
32441=>X"00",
32442=>X"00",
32443=>X"00",
32444=>X"00",
32445=>X"00",
32446=>X"00",
32447=>X"00",
32448=>X"00",
32449=>X"00",
32450=>X"00",
32451=>X"00",
32452=>X"00",
32453=>X"00",
32454=>X"00",
32455=>X"00",
32456=>X"00",
32457=>X"00",
32458=>X"00",
32459=>X"00",
32460=>X"00",
32461=>X"00",
32462=>X"00",
32463=>X"00",
32464=>X"00",
32465=>X"00",
32466=>X"00",
32467=>X"00",
32468=>X"00",
32469=>X"00",
32470=>X"00",
32471=>X"00",
32472=>X"00",
32473=>X"00",
32474=>X"00",
32475=>X"00",
32476=>X"00",
32477=>X"00",
32478=>X"00",
32479=>X"00",
32480=>X"00",
32481=>X"00",
32482=>X"00",
32483=>X"00",
32484=>X"00",
32485=>X"00",
32486=>X"00",
32487=>X"00",
32488=>X"00",
32489=>X"00",
32490=>X"00",
32491=>X"00",
32492=>X"00",
32493=>X"00",
32494=>X"00",
32495=>X"00",
32496=>X"00",
32497=>X"00",
32498=>X"00",
32499=>X"00",
32500=>X"00",
32501=>X"00",
32502=>X"00",
32503=>X"00",
32504=>X"00",
32505=>X"00",
32506=>X"00",
32507=>X"00",
32508=>X"00",
32509=>X"00",
32510=>X"00",
32511=>X"00",
32512=>X"00",
32513=>X"00",
32514=>X"00",
32515=>X"00",
32516=>X"00",
32517=>X"00",
32518=>X"00",
32519=>X"00",
32520=>X"00",
32521=>X"00",
32522=>X"00",
32523=>X"00",
32524=>X"00",
32525=>X"00",
32526=>X"00",
32527=>X"00",
32528=>X"00",
32529=>X"00",
32530=>X"00",
32531=>X"00",
32532=>X"00",
32533=>X"00",
32534=>X"00",
32535=>X"00",
32536=>X"00",
32537=>X"00",
32538=>X"00",
32539=>X"00",
32540=>X"00",
32541=>X"00",
32542=>X"00",
32543=>X"00",
32544=>X"00",
32545=>X"00",
32546=>X"00",
32547=>X"00",
32548=>X"00",
32549=>X"00",
32550=>X"00",
32551=>X"00",
32552=>X"00",
32553=>X"00",
32554=>X"00",
32555=>X"00",
32556=>X"00",
32557=>X"00",
32558=>X"00",
32559=>X"00",
32560=>X"00",
32561=>X"00",
32562=>X"00",
32563=>X"00",
32564=>X"00",
32565=>X"00",
32566=>X"00",
32567=>X"00",
32568=>X"00",
32569=>X"00",
32570=>X"00",
32571=>X"00",
32572=>X"00",
32573=>X"00",
32574=>X"00",
32575=>X"00",
32576=>X"00",
32577=>X"00",
32578=>X"00",
32579=>X"00",
32580=>X"00",
32581=>X"00",
32582=>X"00",
32583=>X"00",
32584=>X"00",
32585=>X"00",
32586=>X"00",
32587=>X"00",
32588=>X"00",
32589=>X"00",
32590=>X"00",
32591=>X"00",
32592=>X"00",
32593=>X"00",
32594=>X"00",
32595=>X"00",
32596=>X"00",
32597=>X"00",
32598=>X"00",
32599=>X"00",
32600=>X"00",
32601=>X"00",
32602=>X"00",
32603=>X"00",
32604=>X"00",
32605=>X"00",
32606=>X"00",
32607=>X"00",
32608=>X"00",
32609=>X"00",
32610=>X"00",
32611=>X"00",
32612=>X"00",
32613=>X"00",
32614=>X"00",
32615=>X"00",
32616=>X"00",
32617=>X"00",
32618=>X"00",
32619=>X"00",
32620=>X"00",
32621=>X"00",
32622=>X"00",
32623=>X"00",
32624=>X"00",
32625=>X"00",
32626=>X"00",
32627=>X"00",
32628=>X"00",
32629=>X"00",
32630=>X"00",
32631=>X"00",
32632=>X"00",
32633=>X"00",
32634=>X"00",
32635=>X"00",
32636=>X"00",
32637=>X"00",
32638=>X"00",
32639=>X"00",
32640=>X"00",
32641=>X"00",
32642=>X"00",
32643=>X"00",
32644=>X"00",
32645=>X"00",
32646=>X"00",
32647=>X"00",
32648=>X"00",
32649=>X"00",
32650=>X"00",
32651=>X"00",
32652=>X"00",
32653=>X"00",
32654=>X"00",
32655=>X"00",
32656=>X"00",
32657=>X"00",
32658=>X"00",
32659=>X"00",
32660=>X"00",
32661=>X"00",
32662=>X"00",
32663=>X"00",
32664=>X"00",
32665=>X"00",
32666=>X"00",
32667=>X"00",
32668=>X"00",
32669=>X"00",
32670=>X"00",
32671=>X"00",
32672=>X"00",
32673=>X"00",
32674=>X"00",
32675=>X"00",
32676=>X"00",
32677=>X"00",
32678=>X"00",
32679=>X"00",
32680=>X"00",
32681=>X"00",
32682=>X"00",
32683=>X"00",
32684=>X"00",
32685=>X"00",
32686=>X"00",
32687=>X"00",
32688=>X"00",
32689=>X"00",
32690=>X"00",
32691=>X"00",
32692=>X"00",
32693=>X"00",
32694=>X"00",
32695=>X"00",
32696=>X"00",
32697=>X"00",
32698=>X"00",
32699=>X"00",
32700=>X"00",
32701=>X"00",
32702=>X"00",
32703=>X"00",
32704=>X"00",
32705=>X"00",
32706=>X"00",
32707=>X"00",
32708=>X"00",
32709=>X"00",
32710=>X"00",
32711=>X"00",
32712=>X"00",
32713=>X"00",
32714=>X"00",
32715=>X"00",
32716=>X"00",
32717=>X"00",
32718=>X"00",
32719=>X"00",
32720=>X"00",
32721=>X"00",
32722=>X"00",
32723=>X"00",
32724=>X"00",
32725=>X"00",
32726=>X"00",
32727=>X"00",
32728=>X"00",
32729=>X"00",
32730=>X"00",
32731=>X"00",
32732=>X"00",
32733=>X"00",
32734=>X"00",
32735=>X"00",
32736=>X"00",
32737=>X"00",
32738=>X"00",
32739=>X"00",
32740=>X"00",
32741=>X"00",
32742=>X"00",
32743=>X"00",
32744=>X"00",
32745=>X"00",
32746=>X"00",
32747=>X"00",
32748=>X"00",
32749=>X"00",
32750=>X"00",
32751=>X"00",
32752=>X"00",
32753=>X"00",
32754=>X"00",
32755=>X"00",
32756=>X"00",
32757=>X"00",
32758=>X"00",
32759=>X"00",
32760=>X"00",
32761=>X"00",
32762=>X"00",
32763=>X"00",
32764=>X"00",
32765=>X"00",
32766=>X"00",
32767=>X"00",
32768=>X"00",
32769=>X"00",
32770=>X"00",
32771=>X"00",
32772=>X"00",
32773=>X"00",
32774=>X"00",
32775=>X"00",
32776=>X"00",
32777=>X"00",
32778=>X"00",
32779=>X"00",
32780=>X"00",
32781=>X"00",
32782=>X"00",
32783=>X"00",
32784=>X"00",
32785=>X"00",
32786=>X"00",
32787=>X"00",
32788=>X"00",
32789=>X"00",
32790=>X"00",
32791=>X"00",
32792=>X"00",
32793=>X"00",
32794=>X"00",
32795=>X"00",
32796=>X"00",
32797=>X"00",
32798=>X"00",
32799=>X"00",
32800=>X"00",
32801=>X"00",
32802=>X"00",
32803=>X"00",
32804=>X"00",
32805=>X"00",
32806=>X"00",
32807=>X"00",
32808=>X"00",
32809=>X"00",
32810=>X"00",
32811=>X"00",
32812=>X"00",
32813=>X"00",
32814=>X"00",
32815=>X"00",
32816=>X"00",
32817=>X"00",
32818=>X"00",
32819=>X"00",
32820=>X"00",
32821=>X"00",
32822=>X"00",
32823=>X"00",
32824=>X"00",
32825=>X"00",
32826=>X"00",
32827=>X"00",
32828=>X"00",
32829=>X"00",
32830=>X"00",
32831=>X"00",
32832=>X"00",
32833=>X"00",
32834=>X"00",
32835=>X"00",
32836=>X"00",
32837=>X"00",
32838=>X"00",
32839=>X"00",
32840=>X"00",
32841=>X"00",
32842=>X"00",
32843=>X"00",
32844=>X"00",
32845=>X"00",
32846=>X"00",
32847=>X"00",
32848=>X"00",
32849=>X"00",
32850=>X"00",
32851=>X"00",
32852=>X"00",
32853=>X"00",
32854=>X"00",
32855=>X"00",
32856=>X"00",
32857=>X"00",
32858=>X"00",
32859=>X"00",
32860=>X"00",
32861=>X"00",
32862=>X"00",
32863=>X"00",
32864=>X"00",
32865=>X"00",
32866=>X"00",
32867=>X"00",
32868=>X"00",
32869=>X"00",
32870=>X"00",
32871=>X"00",
32872=>X"00",
32873=>X"00",
32874=>X"00",
32875=>X"00",
32876=>X"00",
32877=>X"00",
32878=>X"00",
32879=>X"00",
32880=>X"00",
32881=>X"00",
32882=>X"00",
32883=>X"00",
32884=>X"00",
32885=>X"00",
32886=>X"00",
32887=>X"00",
32888=>X"00",
32889=>X"00",
32890=>X"00",
32891=>X"00",
32892=>X"00",
32893=>X"00",
32894=>X"00",
32895=>X"00",
32896=>X"00",
32897=>X"00",
32898=>X"00",
32899=>X"00",
32900=>X"00",
32901=>X"00",
32902=>X"00",
32903=>X"00",
32904=>X"00",
32905=>X"00",
32906=>X"00",
32907=>X"00",
32908=>X"00",
32909=>X"00",
32910=>X"00",
32911=>X"00",
32912=>X"00",
32913=>X"00",
32914=>X"00",
32915=>X"00",
32916=>X"00",
32917=>X"00",
32918=>X"00",
32919=>X"00",
32920=>X"00",
32921=>X"00",
32922=>X"00",
32923=>X"00",
32924=>X"00",
32925=>X"00",
32926=>X"00",
32927=>X"00",
32928=>X"00",
32929=>X"00",
32930=>X"00",
32931=>X"00",
32932=>X"00",
32933=>X"00",
32934=>X"00",
32935=>X"00",
32936=>X"00",
32937=>X"00",
32938=>X"00",
32939=>X"00",
32940=>X"00",
32941=>X"00",
32942=>X"00",
32943=>X"00",
32944=>X"00",
32945=>X"00",
32946=>X"00",
32947=>X"00",
32948=>X"00",
32949=>X"00",
32950=>X"00",
32951=>X"00",
32952=>X"00",
32953=>X"00",
32954=>X"00",
32955=>X"00",
32956=>X"00",
32957=>X"00",
32958=>X"00",
32959=>X"00",
32960=>X"00",
32961=>X"00",
32962=>X"00",
32963=>X"00",
32964=>X"00",
32965=>X"00",
32966=>X"00",
32967=>X"00",
32968=>X"00",
32969=>X"00",
32970=>X"00",
32971=>X"00",
32972=>X"00",
32973=>X"00",
32974=>X"00",
32975=>X"00",
32976=>X"00",
32977=>X"00",
32978=>X"00",
32979=>X"00",
32980=>X"00",
32981=>X"00",
32982=>X"00",
32983=>X"00",
32984=>X"00",
32985=>X"00",
32986=>X"00",
32987=>X"00",
32988=>X"00",
32989=>X"00",
32990=>X"00",
32991=>X"00",
32992=>X"00",
32993=>X"00",
32994=>X"00",
32995=>X"00",
32996=>X"00",
32997=>X"00",
32998=>X"00",
32999=>X"00",
33000=>X"00",
33001=>X"00",
33002=>X"00",
33003=>X"00",
33004=>X"00",
33005=>X"00",
33006=>X"00",
33007=>X"00",
33008=>X"00",
33009=>X"00",
33010=>X"00",
33011=>X"00",
33012=>X"00",
33013=>X"00",
33014=>X"00",
33015=>X"00",
33016=>X"00",
33017=>X"00",
33018=>X"00",
33019=>X"00",
33020=>X"00",
33021=>X"00",
33022=>X"00",
33023=>X"00",
33024=>X"00",
33025=>X"00",
33026=>X"00",
33027=>X"00",
33028=>X"00",
33029=>X"00",
33030=>X"00",
33031=>X"00",
33032=>X"00",
33033=>X"00",
33034=>X"00",
33035=>X"00",
33036=>X"00",
33037=>X"00",
33038=>X"00",
33039=>X"00",
33040=>X"00",
33041=>X"00",
33042=>X"00",
33043=>X"00",
33044=>X"00",
33045=>X"00",
33046=>X"00",
33047=>X"00",
33048=>X"00",
33049=>X"00",
33050=>X"00",
33051=>X"00",
33052=>X"00",
33053=>X"00",
33054=>X"00",
33055=>X"00",
33056=>X"00",
33057=>X"00",
33058=>X"00",
33059=>X"00",
33060=>X"00",
33061=>X"00",
33062=>X"00",
33063=>X"00",
33064=>X"00",
33065=>X"00",
33066=>X"00",
33067=>X"00",
33068=>X"00",
33069=>X"00",
33070=>X"00",
33071=>X"00",
33072=>X"00",
33073=>X"00",
33074=>X"00",
33075=>X"00",
33076=>X"00",
33077=>X"00",
33078=>X"00",
33079=>X"00",
33080=>X"00",
33081=>X"00",
33082=>X"00",
33083=>X"00",
33084=>X"00",
33085=>X"00",
33086=>X"00",
33087=>X"00",
33088=>X"00",
33089=>X"00",
33090=>X"00",
33091=>X"00",
33092=>X"00",
33093=>X"00",
33094=>X"00",
33095=>X"00",
33096=>X"00",
33097=>X"00",
33098=>X"00",
33099=>X"00",
33100=>X"00",
33101=>X"00",
33102=>X"00",
33103=>X"00",
33104=>X"00",
33105=>X"00",
33106=>X"00",
33107=>X"00",
33108=>X"00",
33109=>X"00",
33110=>X"00",
33111=>X"00",
33112=>X"00",
33113=>X"00",
33114=>X"00",
33115=>X"00",
33116=>X"00",
33117=>X"00",
33118=>X"00",
33119=>X"00",
33120=>X"00",
33121=>X"00",
33122=>X"00",
33123=>X"00",
33124=>X"00",
33125=>X"00",
33126=>X"00",
33127=>X"00",
33128=>X"00",
33129=>X"00",
33130=>X"00",
33131=>X"00",
33132=>X"00",
33133=>X"00",
33134=>X"00",
33135=>X"00",
33136=>X"00",
33137=>X"00",
33138=>X"00",
33139=>X"00",
33140=>X"00",
33141=>X"00",
33142=>X"00",
33143=>X"00",
33144=>X"00",
33145=>X"00",
33146=>X"00",
33147=>X"00",
33148=>X"00",
33149=>X"00",
33150=>X"00",
33151=>X"00",
33152=>X"00",
33153=>X"00",
33154=>X"00",
33155=>X"00",
33156=>X"00",
33157=>X"00",
33158=>X"00",
33159=>X"00",
33160=>X"00",
33161=>X"00",
33162=>X"00",
33163=>X"00",
33164=>X"00",
33165=>X"00",
33166=>X"00",
33167=>X"00",
33168=>X"00",
33169=>X"00",
33170=>X"00",
33171=>X"00",
33172=>X"00",
33173=>X"00",
33174=>X"00",
33175=>X"00",
33176=>X"00",
33177=>X"00",
33178=>X"00",
33179=>X"00",
33180=>X"00",
33181=>X"00",
33182=>X"00",
33183=>X"00",
33184=>X"00",
33185=>X"00",
33186=>X"00",
33187=>X"00",
33188=>X"00",
33189=>X"00",
33190=>X"00",
33191=>X"00",
33192=>X"00",
33193=>X"00",
33194=>X"00",
33195=>X"00",
33196=>X"00",
33197=>X"00",
33198=>X"00",
33199=>X"00",
33200=>X"00",
33201=>X"00",
33202=>X"00",
33203=>X"00",
33204=>X"00",
33205=>X"00",
33206=>X"00",
33207=>X"00",
33208=>X"00",
33209=>X"00",
33210=>X"00",
33211=>X"00",
33212=>X"00",
33213=>X"00",
33214=>X"00",
33215=>X"00",
33216=>X"00",
33217=>X"00",
33218=>X"00",
33219=>X"00",
33220=>X"00",
33221=>X"00",
33222=>X"00",
33223=>X"00",
33224=>X"00",
33225=>X"00",
33226=>X"00",
33227=>X"00",
33228=>X"00",
33229=>X"00",
33230=>X"00",
33231=>X"00",
33232=>X"00",
33233=>X"00",
33234=>X"00",
33235=>X"00",
33236=>X"00",
33237=>X"00",
33238=>X"00",
33239=>X"00",
33240=>X"00",
33241=>X"00",
33242=>X"00",
33243=>X"00",
33244=>X"00",
33245=>X"00",
33246=>X"00",
33247=>X"00",
33248=>X"00",
33249=>X"00",
33250=>X"00",
33251=>X"00",
33252=>X"00",
33253=>X"00",
33254=>X"00",
33255=>X"00",
33256=>X"00",
33257=>X"00",
33258=>X"00",
33259=>X"00",
33260=>X"00",
33261=>X"00",
33262=>X"00",
33263=>X"00",
33264=>X"00",
33265=>X"00",
33266=>X"00",
33267=>X"00",
33268=>X"00",
33269=>X"00",
33270=>X"00",
33271=>X"00",
33272=>X"00",
33273=>X"00",
33274=>X"00",
33275=>X"00",
33276=>X"00",
33277=>X"00",
33278=>X"00",
33279=>X"00",
33280=>X"00",
33281=>X"00",
33282=>X"00",
33283=>X"00",
33284=>X"00",
33285=>X"00",
33286=>X"00",
33287=>X"00",
33288=>X"00",
33289=>X"00",
33290=>X"00",
33291=>X"00",
33292=>X"00",
33293=>X"00",
33294=>X"00",
33295=>X"00",
33296=>X"00",
33297=>X"00",
33298=>X"00",
33299=>X"00",
33300=>X"00",
33301=>X"00",
33302=>X"00",
33303=>X"00",
33304=>X"00",
33305=>X"00",
33306=>X"00",
33307=>X"00",
33308=>X"00",
33309=>X"00",
33310=>X"00",
33311=>X"00",
33312=>X"00",
33313=>X"00",
33314=>X"00",
33315=>X"00",
33316=>X"00",
33317=>X"00",
33318=>X"00",
33319=>X"00",
33320=>X"00",
33321=>X"00",
33322=>X"00",
33323=>X"00",
33324=>X"00",
33325=>X"00",
33326=>X"00",
33327=>X"00",
33328=>X"00",
33329=>X"00",
33330=>X"00",
33331=>X"00",
33332=>X"00",
33333=>X"00",
33334=>X"00",
33335=>X"00",
33336=>X"00",
33337=>X"00",
33338=>X"00",
33339=>X"00",
33340=>X"00",
33341=>X"00",
33342=>X"00",
33343=>X"00",
33344=>X"00",
33345=>X"00",
33346=>X"00",
33347=>X"00",
33348=>X"00",
33349=>X"00",
33350=>X"00",
33351=>X"00",
33352=>X"00",
33353=>X"00",
33354=>X"00",
33355=>X"00",
33356=>X"00",
33357=>X"00",
33358=>X"00",
33359=>X"00",
33360=>X"00",
33361=>X"00",
33362=>X"00",
33363=>X"00",
33364=>X"00",
33365=>X"00",
33366=>X"00",
33367=>X"00",
33368=>X"00",
33369=>X"00",
33370=>X"00",
33371=>X"00",
33372=>X"00",
33373=>X"00",
33374=>X"00",
33375=>X"00",
33376=>X"00",
33377=>X"00",
33378=>X"00",
33379=>X"00",
33380=>X"00",
33381=>X"00",
33382=>X"00",
33383=>X"00",
33384=>X"00",
33385=>X"00",
33386=>X"00",
33387=>X"00",
33388=>X"00",
33389=>X"00",
33390=>X"00",
33391=>X"00",
33392=>X"00",
33393=>X"00",
33394=>X"00",
33395=>X"00",
33396=>X"00",
33397=>X"00",
33398=>X"00",
33399=>X"00",
33400=>X"00",
33401=>X"00",
33402=>X"00",
33403=>X"00",
33404=>X"00",
33405=>X"00",
33406=>X"00",
33407=>X"00",
33408=>X"00",
33409=>X"00",
33410=>X"00",
33411=>X"00",
33412=>X"00",
33413=>X"00",
33414=>X"00",
33415=>X"00",
33416=>X"00",
33417=>X"00",
33418=>X"00",
33419=>X"00",
33420=>X"00",
33421=>X"00",
33422=>X"00",
33423=>X"00",
33424=>X"00",
33425=>X"00",
33426=>X"00",
33427=>X"00",
33428=>X"00",
33429=>X"00",
33430=>X"00",
33431=>X"00",
33432=>X"00",
33433=>X"00",
33434=>X"00",
33435=>X"00",
33436=>X"00",
33437=>X"00",
33438=>X"00",
33439=>X"00",
33440=>X"00",
33441=>X"00",
33442=>X"00",
33443=>X"00",
33444=>X"00",
33445=>X"00",
33446=>X"00",
33447=>X"00",
33448=>X"00",
33449=>X"00",
33450=>X"00",
33451=>X"00",
33452=>X"00",
33453=>X"00",
33454=>X"00",
33455=>X"00",
33456=>X"00",
33457=>X"00",
33458=>X"00",
33459=>X"00",
33460=>X"00",
33461=>X"00",
33462=>X"00",
33463=>X"00",
33464=>X"00",
33465=>X"00",
33466=>X"00",
33467=>X"00",
33468=>X"00",
33469=>X"00",
33470=>X"00",
33471=>X"00",
33472=>X"00",
33473=>X"00",
33474=>X"00",
33475=>X"00",
33476=>X"00",
33477=>X"00",
33478=>X"00",
33479=>X"00",
33480=>X"00",
33481=>X"00",
33482=>X"00",
33483=>X"00",
33484=>X"00",
33485=>X"00",
33486=>X"00",
33487=>X"00",
33488=>X"00",
33489=>X"00",
33490=>X"00",
33491=>X"00",
33492=>X"00",
33493=>X"00",
33494=>X"00",
33495=>X"00",
33496=>X"00",
33497=>X"00",
33498=>X"00",
33499=>X"00",
33500=>X"00",
33501=>X"00",
33502=>X"00",
33503=>X"00",
33504=>X"00",
33505=>X"00",
33506=>X"00",
33507=>X"00",
33508=>X"00",
33509=>X"00",
33510=>X"00",
33511=>X"00",
33512=>X"00",
33513=>X"00",
33514=>X"00",
33515=>X"00",
33516=>X"00",
33517=>X"00",
33518=>X"00",
33519=>X"00",
33520=>X"00",
33521=>X"00",
33522=>X"00",
33523=>X"00",
33524=>X"00",
33525=>X"00",
33526=>X"00",
33527=>X"00",
33528=>X"00",
33529=>X"00",
33530=>X"00",
33531=>X"00",
33532=>X"00",
33533=>X"00",
33534=>X"00",
33535=>X"00",
33536=>X"00",
33537=>X"00",
33538=>X"00",
33539=>X"00",
33540=>X"00",
33541=>X"00",
33542=>X"00",
33543=>X"00",
33544=>X"00",
33545=>X"00",
33546=>X"00",
33547=>X"00",
33548=>X"00",
33549=>X"00",
33550=>X"00",
33551=>X"00",
33552=>X"00",
33553=>X"00",
33554=>X"00",
33555=>X"00",
33556=>X"00",
33557=>X"00",
33558=>X"00",
33559=>X"00",
33560=>X"00",
33561=>X"00",
33562=>X"00",
33563=>X"00",
33564=>X"00",
33565=>X"00",
33566=>X"00",
33567=>X"00",
33568=>X"00",
33569=>X"00",
33570=>X"00",
33571=>X"00",
33572=>X"00",
33573=>X"00",
33574=>X"00",
33575=>X"00",
33576=>X"00",
33577=>X"00",
33578=>X"00",
33579=>X"00",
33580=>X"00",
33581=>X"00",
33582=>X"00",
33583=>X"00",
33584=>X"00",
33585=>X"00",
33586=>X"00",
33587=>X"00",
33588=>X"00",
33589=>X"00",
33590=>X"00",
33591=>X"00",
33592=>X"00",
33593=>X"00",
33594=>X"00",
33595=>X"00",
33596=>X"00",
33597=>X"00",
33598=>X"00",
33599=>X"00",
33600=>X"00",
33601=>X"00",
33602=>X"00",
33603=>X"00",
33604=>X"00",
33605=>X"00",
33606=>X"00",
33607=>X"00",
33608=>X"00",
33609=>X"00",
33610=>X"00",
33611=>X"00",
33612=>X"00",
33613=>X"00",
33614=>X"00",
33615=>X"00",
33616=>X"00",
33617=>X"00",
33618=>X"00",
33619=>X"00",
33620=>X"00",
33621=>X"00",
33622=>X"00",
33623=>X"00",
33624=>X"00",
33625=>X"00",
33626=>X"00",
33627=>X"00",
33628=>X"00",
33629=>X"00",
33630=>X"00",
33631=>X"00",
33632=>X"00",
33633=>X"00",
33634=>X"00",
33635=>X"00",
33636=>X"00",
33637=>X"00",
33638=>X"00",
33639=>X"00",
33640=>X"00",
33641=>X"00",
33642=>X"00",
33643=>X"00",
33644=>X"00",
33645=>X"00",
33646=>X"00",
33647=>X"00",
33648=>X"00",
33649=>X"00",
33650=>X"00",
33651=>X"00",
33652=>X"00",
33653=>X"00",
33654=>X"00",
33655=>X"00",
33656=>X"00",
33657=>X"00",
33658=>X"00",
33659=>X"00",
33660=>X"00",
33661=>X"00",
33662=>X"00",
33663=>X"00",
33664=>X"00",
33665=>X"00",
33666=>X"00",
33667=>X"00",
33668=>X"00",
33669=>X"00",
33670=>X"00",
33671=>X"00",
33672=>X"00",
33673=>X"00",
33674=>X"00",
33675=>X"00",
33676=>X"00",
33677=>X"00",
33678=>X"00",
33679=>X"00",
33680=>X"00",
33681=>X"00",
33682=>X"00",
33683=>X"00",
33684=>X"00",
33685=>X"00",
33686=>X"00",
33687=>X"00",
33688=>X"00",
33689=>X"00",
33690=>X"00",
33691=>X"00",
33692=>X"00",
33693=>X"00",
33694=>X"00",
33695=>X"00",
33696=>X"00",
33697=>X"00",
33698=>X"00",
33699=>X"00",
33700=>X"00",
33701=>X"00",
33702=>X"00",
33703=>X"00",
33704=>X"00",
33705=>X"00",
33706=>X"00",
33707=>X"00",
33708=>X"00",
33709=>X"00",
33710=>X"00",
33711=>X"00",
33712=>X"00",
33713=>X"00",
33714=>X"00",
33715=>X"00",
33716=>X"00",
33717=>X"00",
33718=>X"00",
33719=>X"00",
33720=>X"00",
33721=>X"00",
33722=>X"00",
33723=>X"00",
33724=>X"00",
33725=>X"00",
33726=>X"00",
33727=>X"00",
33728=>X"00",
33729=>X"00",
33730=>X"00",
33731=>X"00",
33732=>X"00",
33733=>X"00",
33734=>X"00",
33735=>X"00",
33736=>X"00",
33737=>X"00",
33738=>X"00",
33739=>X"00",
33740=>X"00",
33741=>X"00",
33742=>X"00",
33743=>X"00",
33744=>X"00",
33745=>X"00",
33746=>X"00",
33747=>X"00",
33748=>X"00",
33749=>X"00",
33750=>X"00",
33751=>X"00",
33752=>X"00",
33753=>X"00",
33754=>X"00",
33755=>X"00",
33756=>X"00",
33757=>X"00",
33758=>X"00",
33759=>X"00",
33760=>X"00",
33761=>X"00",
33762=>X"00",
33763=>X"00",
33764=>X"00",
33765=>X"00",
33766=>X"00",
33767=>X"00",
33768=>X"00",
33769=>X"00",
33770=>X"00",
33771=>X"00",
33772=>X"00",
33773=>X"00",
33774=>X"00",
33775=>X"00",
33776=>X"00",
33777=>X"00",
33778=>X"00",
33779=>X"00",
33780=>X"00",
33781=>X"00",
33782=>X"00",
33783=>X"00",
33784=>X"00",
33785=>X"00",
33786=>X"00",
33787=>X"00",
33788=>X"00",
33789=>X"00",
33790=>X"00",
33791=>X"00",
33792=>X"00",
33793=>X"00",
33794=>X"00",
33795=>X"00",
33796=>X"00",
33797=>X"00",
33798=>X"00",
33799=>X"00",
33800=>X"00",
33801=>X"00",
33802=>X"00",
33803=>X"00",
33804=>X"00",
33805=>X"00",
33806=>X"00",
33807=>X"00",
33808=>X"00",
33809=>X"00",
33810=>X"00",
33811=>X"00",
33812=>X"00",
33813=>X"00",
33814=>X"00",
33815=>X"00",
33816=>X"00",
33817=>X"00",
33818=>X"00",
33819=>X"00",
33820=>X"00",
33821=>X"00",
33822=>X"00",
33823=>X"00",
33824=>X"00",
33825=>X"00",
33826=>X"00",
33827=>X"00",
33828=>X"00",
33829=>X"00",
33830=>X"00",
33831=>X"00",
33832=>X"00",
33833=>X"00",
33834=>X"00",
33835=>X"00",
33836=>X"00",
33837=>X"00",
33838=>X"00",
33839=>X"00",
33840=>X"00",
33841=>X"00",
33842=>X"00",
33843=>X"00",
33844=>X"00",
33845=>X"00",
33846=>X"00",
33847=>X"00",
33848=>X"00",
33849=>X"00",
33850=>X"00",
33851=>X"00",
33852=>X"00",
33853=>X"00",
33854=>X"00",
33855=>X"00",
33856=>X"00",
33857=>X"00",
33858=>X"00",
33859=>X"00",
33860=>X"00",
33861=>X"00",
33862=>X"00",
33863=>X"00",
33864=>X"00",
33865=>X"00",
33866=>X"00",
33867=>X"00",
33868=>X"00",
33869=>X"00",
33870=>X"00",
33871=>X"00",
33872=>X"00",
33873=>X"00",
33874=>X"00",
33875=>X"00",
33876=>X"00",
33877=>X"00",
33878=>X"00",
33879=>X"00",
33880=>X"00",
33881=>X"00",
33882=>X"00",
33883=>X"00",
33884=>X"00",
33885=>X"00",
33886=>X"00",
33887=>X"00",
33888=>X"00",
33889=>X"00",
33890=>X"00",
33891=>X"00",
33892=>X"00",
33893=>X"00",
33894=>X"00",
33895=>X"00",
33896=>X"00",
33897=>X"00",
33898=>X"00",
33899=>X"00",
33900=>X"00",
33901=>X"00",
33902=>X"00",
33903=>X"00",
33904=>X"00",
33905=>X"00",
33906=>X"00",
33907=>X"00",
33908=>X"00",
33909=>X"00",
33910=>X"00",
33911=>X"00",
33912=>X"00",
33913=>X"00",
33914=>X"00",
33915=>X"00",
33916=>X"00",
33917=>X"00",
33918=>X"00",
33919=>X"00",
33920=>X"00",
33921=>X"00",
33922=>X"00",
33923=>X"00",
33924=>X"00",
33925=>X"00",
33926=>X"00",
33927=>X"00",
33928=>X"00",
33929=>X"00",
33930=>X"00",
33931=>X"00",
33932=>X"00",
33933=>X"00",
33934=>X"00",
33935=>X"00",
33936=>X"00",
33937=>X"00",
33938=>X"00",
33939=>X"00",
33940=>X"00",
33941=>X"00",
33942=>X"00",
33943=>X"00",
33944=>X"00",
33945=>X"00",
33946=>X"00",
33947=>X"00",
33948=>X"00",
33949=>X"00",
33950=>X"00",
33951=>X"00",
33952=>X"00",
33953=>X"00",
33954=>X"00",
33955=>X"00",
33956=>X"00",
33957=>X"00",
33958=>X"00",
33959=>X"00",
33960=>X"00",
33961=>X"00",
33962=>X"00",
33963=>X"00",
33964=>X"00",
33965=>X"00",
33966=>X"00",
33967=>X"00",
33968=>X"00",
33969=>X"00",
33970=>X"00",
33971=>X"00",
33972=>X"00",
33973=>X"00",
33974=>X"00",
33975=>X"00",
33976=>X"00",
33977=>X"00",
33978=>X"00",
33979=>X"00",
33980=>X"00",
33981=>X"00",
33982=>X"00",
33983=>X"00",
33984=>X"00",
33985=>X"00",
33986=>X"00",
33987=>X"00",
33988=>X"00",
33989=>X"00",
33990=>X"00",
33991=>X"00",
33992=>X"00",
33993=>X"00",
33994=>X"00",
33995=>X"00",
33996=>X"00",
33997=>X"00",
33998=>X"00",
33999=>X"00",
34000=>X"00",
34001=>X"00",
34002=>X"00",
34003=>X"00",
34004=>X"00",
34005=>X"00",
34006=>X"00",
34007=>X"00",
34008=>X"00",
34009=>X"00",
34010=>X"00",
34011=>X"00",
34012=>X"00",
34013=>X"00",
34014=>X"00",
34015=>X"00",
34016=>X"00",
34017=>X"00",
34018=>X"00",
34019=>X"00",
34020=>X"00",
34021=>X"00",
34022=>X"00",
34023=>X"00",
34024=>X"00",
34025=>X"00",
34026=>X"00",
34027=>X"00",
34028=>X"00",
34029=>X"00",
34030=>X"00",
34031=>X"00",
34032=>X"00",
34033=>X"00",
34034=>X"00",
34035=>X"00",
34036=>X"00",
34037=>X"00",
34038=>X"00",
34039=>X"00",
34040=>X"00",
34041=>X"00",
34042=>X"00",
34043=>X"00",
34044=>X"00",
34045=>X"00",
34046=>X"00",
34047=>X"00",
34048=>X"00",
34049=>X"00",
34050=>X"00",
34051=>X"00",
34052=>X"00",
34053=>X"00",
34054=>X"00",
34055=>X"00",
34056=>X"00",
34057=>X"00",
34058=>X"00",
34059=>X"00",
34060=>X"00",
34061=>X"00",
34062=>X"00",
34063=>X"00",
34064=>X"00",
34065=>X"00",
34066=>X"00",
34067=>X"00",
34068=>X"00",
34069=>X"00",
34070=>X"00",
34071=>X"00",
34072=>X"00",
34073=>X"00",
34074=>X"00",
34075=>X"00",
34076=>X"00",
34077=>X"00",
34078=>X"00",
34079=>X"00",
34080=>X"00",
34081=>X"00",
34082=>X"00",
34083=>X"00",
34084=>X"00",
34085=>X"00",
34086=>X"00",
34087=>X"00",
34088=>X"00",
34089=>X"00",
34090=>X"00",
34091=>X"00",
34092=>X"00",
34093=>X"00",
34094=>X"00",
34095=>X"00",
34096=>X"00",
34097=>X"00",
34098=>X"00",
34099=>X"00",
34100=>X"00",
34101=>X"00",
34102=>X"00",
34103=>X"00",
34104=>X"00",
34105=>X"00",
34106=>X"00",
34107=>X"00",
34108=>X"00",
34109=>X"00",
34110=>X"00",
34111=>X"00",
34112=>X"00",
34113=>X"00",
34114=>X"00",
34115=>X"00",
34116=>X"00",
34117=>X"00",
34118=>X"00",
34119=>X"00",
34120=>X"00",
34121=>X"00",
34122=>X"00",
34123=>X"00",
34124=>X"00",
34125=>X"00",
34126=>X"00",
34127=>X"00",
34128=>X"00",
34129=>X"00",
34130=>X"00",
34131=>X"00",
34132=>X"00",
34133=>X"00",
34134=>X"00",
34135=>X"00",
34136=>X"00",
34137=>X"00",
34138=>X"00",
34139=>X"00",
34140=>X"00",
34141=>X"00",
34142=>X"00",
34143=>X"00",
34144=>X"00",
34145=>X"00",
34146=>X"00",
34147=>X"00",
34148=>X"00",
34149=>X"00",
34150=>X"00",
34151=>X"00",
34152=>X"00",
34153=>X"00",
34154=>X"00",
34155=>X"00",
34156=>X"00",
34157=>X"00",
34158=>X"00",
34159=>X"00",
34160=>X"00",
34161=>X"00",
34162=>X"00",
34163=>X"00",
34164=>X"00",
34165=>X"00",
34166=>X"00",
34167=>X"00",
34168=>X"00",
34169=>X"00",
34170=>X"00",
34171=>X"00",
34172=>X"00",
34173=>X"00",
34174=>X"00",
34175=>X"00",
34176=>X"00",
34177=>X"00",
34178=>X"00",
34179=>X"00",
34180=>X"00",
34181=>X"00",
34182=>X"00",
34183=>X"00",
34184=>X"00",
34185=>X"00",
34186=>X"00",
34187=>X"00",
34188=>X"00",
34189=>X"00",
34190=>X"00",
34191=>X"00",
34192=>X"00",
34193=>X"00",
34194=>X"00",
34195=>X"00",
34196=>X"00",
34197=>X"00",
34198=>X"00",
34199=>X"00",
34200=>X"00",
34201=>X"00",
34202=>X"00",
34203=>X"00",
34204=>X"00",
34205=>X"00",
34206=>X"00",
34207=>X"00",
34208=>X"00",
34209=>X"00",
34210=>X"00",
34211=>X"00",
34212=>X"00",
34213=>X"00",
34214=>X"00",
34215=>X"00",
34216=>X"00",
34217=>X"00",
34218=>X"00",
34219=>X"00",
34220=>X"00",
34221=>X"00",
34222=>X"00",
34223=>X"00",
34224=>X"00",
34225=>X"00",
34226=>X"00",
34227=>X"00",
34228=>X"00",
34229=>X"00",
34230=>X"00",
34231=>X"00",
34232=>X"00",
34233=>X"00",
34234=>X"00",
34235=>X"00",
34236=>X"00",
34237=>X"00",
34238=>X"00",
34239=>X"00",
34240=>X"00",
34241=>X"00",
34242=>X"00",
34243=>X"00",
34244=>X"00",
34245=>X"00",
34246=>X"00",
34247=>X"00",
34248=>X"00",
34249=>X"00",
34250=>X"00",
34251=>X"00",
34252=>X"00",
34253=>X"00",
34254=>X"00",
34255=>X"00",
34256=>X"00",
34257=>X"00",
34258=>X"00",
34259=>X"00",
34260=>X"00",
34261=>X"00",
34262=>X"00",
34263=>X"00",
34264=>X"00",
34265=>X"00",
34266=>X"00",
34267=>X"00",
34268=>X"00",
34269=>X"00",
34270=>X"00",
34271=>X"00",
34272=>X"00",
34273=>X"00",
34274=>X"00",
34275=>X"00",
34276=>X"00",
34277=>X"00",
34278=>X"00",
34279=>X"00",
34280=>X"00",
34281=>X"00",
34282=>X"00",
34283=>X"00",
34284=>X"00",
34285=>X"00",
34286=>X"00",
34287=>X"00",
34288=>X"00",
34289=>X"00",
34290=>X"00",
34291=>X"00",
34292=>X"00",
34293=>X"00",
34294=>X"00",
34295=>X"00",
34296=>X"00",
34297=>X"00",
34298=>X"00",
34299=>X"00",
34300=>X"00",
34301=>X"00",
34302=>X"00",
34303=>X"00",
34304=>X"00",
34305=>X"00",
34306=>X"00",
34307=>X"00",
34308=>X"00",
34309=>X"00",
34310=>X"00",
34311=>X"00",
34312=>X"00",
34313=>X"00",
34314=>X"00",
34315=>X"00",
34316=>X"00",
34317=>X"00",
34318=>X"00",
34319=>X"00",
34320=>X"00",
34321=>X"00",
34322=>X"00",
34323=>X"00",
34324=>X"00",
34325=>X"00",
34326=>X"00",
34327=>X"00",
34328=>X"00",
34329=>X"00",
34330=>X"00",
34331=>X"00",
34332=>X"00",
34333=>X"00",
34334=>X"00",
34335=>X"00",
34336=>X"00",
34337=>X"00",
34338=>X"00",
34339=>X"00",
34340=>X"00",
34341=>X"00",
34342=>X"00",
34343=>X"00",
34344=>X"00",
34345=>X"00",
34346=>X"00",
34347=>X"00",
34348=>X"00",
34349=>X"00",
34350=>X"00",
34351=>X"00",
34352=>X"00",
34353=>X"00",
34354=>X"00",
34355=>X"00",
34356=>X"00",
34357=>X"00",
34358=>X"00",
34359=>X"00",
34360=>X"00",
34361=>X"00",
34362=>X"00",
34363=>X"00",
34364=>X"00",
34365=>X"00",
34366=>X"00",
34367=>X"00",
34368=>X"00",
34369=>X"00",
34370=>X"00",
34371=>X"00",
34372=>X"00",
34373=>X"00",
34374=>X"00",
34375=>X"00",
34376=>X"00",
34377=>X"00",
34378=>X"00",
34379=>X"00",
34380=>X"00",
34381=>X"00",
34382=>X"00",
34383=>X"00",
34384=>X"00",
34385=>X"00",
34386=>X"00",
34387=>X"00",
34388=>X"00",
34389=>X"00",
34390=>X"00",
34391=>X"00",
34392=>X"00",
34393=>X"00",
34394=>X"00",
34395=>X"00",
34396=>X"00",
34397=>X"00",
34398=>X"00",
34399=>X"00",
34400=>X"00",
34401=>X"00",
34402=>X"00",
34403=>X"00",
34404=>X"00",
34405=>X"00",
34406=>X"00",
34407=>X"00",
34408=>X"00",
34409=>X"00",
34410=>X"00",
34411=>X"00",
34412=>X"00",
34413=>X"00",
34414=>X"00",
34415=>X"00",
34416=>X"00",
34417=>X"00",
34418=>X"00",
34419=>X"00",
34420=>X"00",
34421=>X"00",
34422=>X"00",
34423=>X"00",
34424=>X"00",
34425=>X"00",
34426=>X"00",
34427=>X"00",
34428=>X"00",
34429=>X"00",
34430=>X"00",
34431=>X"00",
34432=>X"00",
34433=>X"00",
34434=>X"00",
34435=>X"00",
34436=>X"00",
34437=>X"00",
34438=>X"00",
34439=>X"00",
34440=>X"00",
34441=>X"00",
34442=>X"00",
34443=>X"00",
34444=>X"00",
34445=>X"00",
34446=>X"00",
34447=>X"00",
34448=>X"00",
34449=>X"00",
34450=>X"00",
34451=>X"00",
34452=>X"00",
34453=>X"00",
34454=>X"00",
34455=>X"00",
34456=>X"00",
34457=>X"00",
34458=>X"00",
34459=>X"00",
34460=>X"00",
34461=>X"00",
34462=>X"00",
34463=>X"00",
34464=>X"00",
34465=>X"00",
34466=>X"00",
34467=>X"00",
34468=>X"00",
34469=>X"00",
34470=>X"00",
34471=>X"00",
34472=>X"00",
34473=>X"00",
34474=>X"00",
34475=>X"00",
34476=>X"00",
34477=>X"00",
34478=>X"00",
34479=>X"00",
34480=>X"00",
34481=>X"00",
34482=>X"00",
34483=>X"00",
34484=>X"00",
34485=>X"00",
34486=>X"00",
34487=>X"00",
34488=>X"00",
34489=>X"00",
34490=>X"00",
34491=>X"00",
34492=>X"00",
34493=>X"00",
34494=>X"00",
34495=>X"00",
34496=>X"00",
34497=>X"00",
34498=>X"00",
34499=>X"00",
34500=>X"00",
34501=>X"00",
34502=>X"00",
34503=>X"00",
34504=>X"00",
34505=>X"00",
34506=>X"00",
34507=>X"00",
34508=>X"00",
34509=>X"00",
34510=>X"00",
34511=>X"00",
34512=>X"00",
34513=>X"00",
34514=>X"00",
34515=>X"00",
34516=>X"00",
34517=>X"00",
34518=>X"00",
34519=>X"00",
34520=>X"00",
34521=>X"00",
34522=>X"00",
34523=>X"00",
34524=>X"00",
34525=>X"00",
34526=>X"00",
34527=>X"00",
34528=>X"00",
34529=>X"00",
34530=>X"00",
34531=>X"00",
34532=>X"00",
34533=>X"00",
34534=>X"00",
34535=>X"00",
34536=>X"00",
34537=>X"00",
34538=>X"00",
34539=>X"00",
34540=>X"00",
34541=>X"00",
34542=>X"00",
34543=>X"00",
34544=>X"00",
34545=>X"00",
34546=>X"00",
34547=>X"00",
34548=>X"00",
34549=>X"00",
34550=>X"00",
34551=>X"00",
34552=>X"00",
34553=>X"00",
34554=>X"00",
34555=>X"00",
34556=>X"00",
34557=>X"00",
34558=>X"00",
34559=>X"00",
34560=>X"00",
34561=>X"00",
34562=>X"00",
34563=>X"00",
34564=>X"00",
34565=>X"00",
34566=>X"00",
34567=>X"00",
34568=>X"00",
34569=>X"00",
34570=>X"00",
34571=>X"00",
34572=>X"00",
34573=>X"00",
34574=>X"00",
34575=>X"00",
34576=>X"00",
34577=>X"00",
34578=>X"00",
34579=>X"00",
34580=>X"00",
34581=>X"00",
34582=>X"00",
34583=>X"00",
34584=>X"00",
34585=>X"00",
34586=>X"00",
34587=>X"00",
34588=>X"00",
34589=>X"00",
34590=>X"00",
34591=>X"00",
34592=>X"00",
34593=>X"00",
34594=>X"00",
34595=>X"00",
34596=>X"00",
34597=>X"00",
34598=>X"00",
34599=>X"00",
34600=>X"00",
34601=>X"00",
34602=>X"00",
34603=>X"00",
34604=>X"00",
34605=>X"00",
34606=>X"00",
34607=>X"00",
34608=>X"00",
34609=>X"00",
34610=>X"00",
34611=>X"00",
34612=>X"00",
34613=>X"00",
34614=>X"00",
34615=>X"00",
34616=>X"00",
34617=>X"00",
34618=>X"00",
34619=>X"00",
34620=>X"00",
34621=>X"00",
34622=>X"00",
34623=>X"00",
34624=>X"00",
34625=>X"00",
34626=>X"00",
34627=>X"00",
34628=>X"00",
34629=>X"00",
34630=>X"00",
34631=>X"00",
34632=>X"00",
34633=>X"00",
34634=>X"00",
34635=>X"00",
34636=>X"00",
34637=>X"00",
34638=>X"00",
34639=>X"00",
34640=>X"00",
34641=>X"00",
34642=>X"00",
34643=>X"00",
34644=>X"00",
34645=>X"00",
34646=>X"00",
34647=>X"00",
34648=>X"00",
34649=>X"00",
34650=>X"00",
34651=>X"00",
34652=>X"00",
34653=>X"00",
34654=>X"00",
34655=>X"00",
34656=>X"00",
34657=>X"00",
34658=>X"00",
34659=>X"00",
34660=>X"00",
34661=>X"00",
34662=>X"00",
34663=>X"00",
34664=>X"00",
34665=>X"00",
34666=>X"00",
34667=>X"00",
34668=>X"00",
34669=>X"00",
34670=>X"00",
34671=>X"00",
34672=>X"00",
34673=>X"00",
34674=>X"00",
34675=>X"00",
34676=>X"00",
34677=>X"00",
34678=>X"00",
34679=>X"00",
34680=>X"00",
34681=>X"00",
34682=>X"00",
34683=>X"00",
34684=>X"00",
34685=>X"00",
34686=>X"00",
34687=>X"00",
34688=>X"00",
34689=>X"00",
34690=>X"00",
34691=>X"00",
34692=>X"00",
34693=>X"00",
34694=>X"00",
34695=>X"00",
34696=>X"00",
34697=>X"00",
34698=>X"00",
34699=>X"00",
34700=>X"00",
34701=>X"00",
34702=>X"00",
34703=>X"00",
34704=>X"00",
34705=>X"00",
34706=>X"00",
34707=>X"00",
34708=>X"00",
34709=>X"00",
34710=>X"00",
34711=>X"00",
34712=>X"00",
34713=>X"00",
34714=>X"00",
34715=>X"00",
34716=>X"00",
34717=>X"00",
34718=>X"00",
34719=>X"00",
34720=>X"00",
34721=>X"00",
34722=>X"00",
34723=>X"00",
34724=>X"00",
34725=>X"00",
34726=>X"00",
34727=>X"00",
34728=>X"00",
34729=>X"00",
34730=>X"00",
34731=>X"00",
34732=>X"00",
34733=>X"00",
34734=>X"00",
34735=>X"00",
34736=>X"00",
34737=>X"00",
34738=>X"00",
34739=>X"00",
34740=>X"00",
34741=>X"00",
34742=>X"00",
34743=>X"00",
34744=>X"00",
34745=>X"00",
34746=>X"00",
34747=>X"00",
34748=>X"00",
34749=>X"00",
34750=>X"00",
34751=>X"00",
34752=>X"00",
34753=>X"00",
34754=>X"00",
34755=>X"00",
34756=>X"00",
34757=>X"00",
34758=>X"00",
34759=>X"00",
34760=>X"00",
34761=>X"00",
34762=>X"00",
34763=>X"00",
34764=>X"00",
34765=>X"00",
34766=>X"00",
34767=>X"00",
34768=>X"00",
34769=>X"00",
34770=>X"00",
34771=>X"00",
34772=>X"00",
34773=>X"00",
34774=>X"00",
34775=>X"00",
34776=>X"00",
34777=>X"00",
34778=>X"00",
34779=>X"00",
34780=>X"00",
34781=>X"00",
34782=>X"00",
34783=>X"00",
34784=>X"00",
34785=>X"00",
34786=>X"00",
34787=>X"00",
34788=>X"00",
34789=>X"00",
34790=>X"00",
34791=>X"00",
34792=>X"00",
34793=>X"00",
34794=>X"00",
34795=>X"00",
34796=>X"00",
34797=>X"00",
34798=>X"00",
34799=>X"00",
34800=>X"00",
34801=>X"00",
34802=>X"00",
34803=>X"00",
34804=>X"00",
34805=>X"00",
34806=>X"00",
34807=>X"00",
34808=>X"00",
34809=>X"00",
34810=>X"00",
34811=>X"00",
34812=>X"00",
34813=>X"00",
34814=>X"00",
34815=>X"00",
34816=>X"00",
34817=>X"00",
34818=>X"00",
34819=>X"00",
34820=>X"00",
34821=>X"00",
34822=>X"00",
34823=>X"00",
34824=>X"00",
34825=>X"00",
34826=>X"00",
34827=>X"00",
34828=>X"00",
34829=>X"00",
34830=>X"00",
34831=>X"00",
34832=>X"00",
34833=>X"00",
34834=>X"00",
34835=>X"00",
34836=>X"00",
34837=>X"00",
34838=>X"00",
34839=>X"00",
34840=>X"00",
34841=>X"00",
34842=>X"00",
34843=>X"00",
34844=>X"00",
34845=>X"00",
34846=>X"00",
34847=>X"00",
34848=>X"00",
34849=>X"00",
34850=>X"00",
34851=>X"00",
34852=>X"00",
34853=>X"00",
34854=>X"00",
34855=>X"00",
34856=>X"00",
34857=>X"00",
34858=>X"00",
34859=>X"00",
34860=>X"00",
34861=>X"00",
34862=>X"00",
34863=>X"00",
34864=>X"00",
34865=>X"00",
34866=>X"00",
34867=>X"00",
34868=>X"00",
34869=>X"00",
34870=>X"00",
34871=>X"00",
34872=>X"00",
34873=>X"00",
34874=>X"00",
34875=>X"00",
34876=>X"00",
34877=>X"00",
34878=>X"00",
34879=>X"00",
34880=>X"00",
34881=>X"00",
34882=>X"00",
34883=>X"00",
34884=>X"00",
34885=>X"00",
34886=>X"00",
34887=>X"00",
34888=>X"00",
34889=>X"00",
34890=>X"00",
34891=>X"00",
34892=>X"00",
34893=>X"00",
34894=>X"00",
34895=>X"00",
34896=>X"00",
34897=>X"00",
34898=>X"00",
34899=>X"00",
34900=>X"00",
34901=>X"00",
34902=>X"00",
34903=>X"00",
34904=>X"00",
34905=>X"00",
34906=>X"00",
34907=>X"00",
34908=>X"00",
34909=>X"00",
34910=>X"00",
34911=>X"00",
34912=>X"00",
34913=>X"00",
34914=>X"00",
34915=>X"00",
34916=>X"00",
34917=>X"00",
34918=>X"00",
34919=>X"00",
34920=>X"00",
34921=>X"00",
34922=>X"00",
34923=>X"00",
34924=>X"00",
34925=>X"00",
34926=>X"00",
34927=>X"00",
34928=>X"00",
34929=>X"00",
34930=>X"00",
34931=>X"00",
34932=>X"00",
34933=>X"00",
34934=>X"00",
34935=>X"00",
34936=>X"00",
34937=>X"00",
34938=>X"00",
34939=>X"00",
34940=>X"00",
34941=>X"00",
34942=>X"00",
34943=>X"00",
34944=>X"00",
34945=>X"00",
34946=>X"00",
34947=>X"00",
34948=>X"00",
34949=>X"00",
34950=>X"00",
34951=>X"00",
34952=>X"00",
34953=>X"00",
34954=>X"00",
34955=>X"00",
34956=>X"00",
34957=>X"00",
34958=>X"00",
34959=>X"00",
34960=>X"00",
34961=>X"00",
34962=>X"00",
34963=>X"00",
34964=>X"00",
34965=>X"00",
34966=>X"00",
34967=>X"00",
34968=>X"00",
34969=>X"00",
34970=>X"00",
34971=>X"00",
34972=>X"00",
34973=>X"00",
34974=>X"00",
34975=>X"00",
34976=>X"00",
34977=>X"00",
34978=>X"00",
34979=>X"00",
34980=>X"00",
34981=>X"00",
34982=>X"00",
34983=>X"00",
34984=>X"00",
34985=>X"00",
34986=>X"00",
34987=>X"00",
34988=>X"00",
34989=>X"00",
34990=>X"00",
34991=>X"00",
34992=>X"00",
34993=>X"00",
34994=>X"00",
34995=>X"00",
34996=>X"00",
34997=>X"00",
34998=>X"00",
34999=>X"00",
35000=>X"00",
35001=>X"00",
35002=>X"00",
35003=>X"00",
35004=>X"00",
35005=>X"00",
35006=>X"00",
35007=>X"00",
35008=>X"00",
35009=>X"00",
35010=>X"00",
35011=>X"00",
35012=>X"00",
35013=>X"00",
35014=>X"00",
35015=>X"00",
35016=>X"00",
35017=>X"00",
35018=>X"00",
35019=>X"00",
35020=>X"00",
35021=>X"00",
35022=>X"00",
35023=>X"00",
35024=>X"00",
35025=>X"00",
35026=>X"00",
35027=>X"00",
35028=>X"00",
35029=>X"00",
35030=>X"00",
35031=>X"00",
35032=>X"00",
35033=>X"00",
35034=>X"00",
35035=>X"00",
35036=>X"00",
35037=>X"00",
35038=>X"00",
35039=>X"00",
35040=>X"00",
35041=>X"00",
35042=>X"00",
35043=>X"00",
35044=>X"00",
35045=>X"00",
35046=>X"00",
35047=>X"00",
35048=>X"00",
35049=>X"00",
35050=>X"00",
35051=>X"00",
35052=>X"00",
35053=>X"00",
35054=>X"00",
35055=>X"00",
35056=>X"00",
35057=>X"00",
35058=>X"00",
35059=>X"00",
35060=>X"00",
35061=>X"00",
35062=>X"00",
35063=>X"00",
35064=>X"00",
35065=>X"00",
35066=>X"00",
35067=>X"00",
35068=>X"00",
35069=>X"00",
35070=>X"00",
35071=>X"00",
35072=>X"00",
35073=>X"00",
35074=>X"00",
35075=>X"00",
35076=>X"00",
35077=>X"00",
35078=>X"00",
35079=>X"00",
35080=>X"00",
35081=>X"00",
35082=>X"00",
35083=>X"00",
35084=>X"00",
35085=>X"00",
35086=>X"00",
35087=>X"00",
35088=>X"00",
35089=>X"00",
35090=>X"00",
35091=>X"00",
35092=>X"00",
35093=>X"00",
35094=>X"00",
35095=>X"00",
35096=>X"00",
35097=>X"00",
35098=>X"00",
35099=>X"00",
35100=>X"00",
35101=>X"00",
35102=>X"00",
35103=>X"00",
35104=>X"00",
35105=>X"00",
35106=>X"00",
35107=>X"00",
35108=>X"00",
35109=>X"00",
35110=>X"00",
35111=>X"00",
35112=>X"00",
35113=>X"00",
35114=>X"00",
35115=>X"00",
35116=>X"00",
35117=>X"00",
35118=>X"00",
35119=>X"00",
35120=>X"00",
35121=>X"00",
35122=>X"00",
35123=>X"00",
35124=>X"00",
35125=>X"00",
35126=>X"00",
35127=>X"00",
35128=>X"00",
35129=>X"00",
35130=>X"00",
35131=>X"00",
35132=>X"00",
35133=>X"00",
35134=>X"00",
35135=>X"00",
35136=>X"00",
35137=>X"00",
35138=>X"00",
35139=>X"00",
35140=>X"00",
35141=>X"00",
35142=>X"00",
35143=>X"00",
35144=>X"00",
35145=>X"00",
35146=>X"00",
35147=>X"00",
35148=>X"00",
35149=>X"00",
35150=>X"00",
35151=>X"00",
35152=>X"00",
35153=>X"00",
35154=>X"00",
35155=>X"00",
35156=>X"00",
35157=>X"00",
35158=>X"00",
35159=>X"00",
35160=>X"00",
35161=>X"00",
35162=>X"00",
35163=>X"00",
35164=>X"00",
35165=>X"00",
35166=>X"00",
35167=>X"00",
35168=>X"00",
35169=>X"00",
35170=>X"00",
35171=>X"00",
35172=>X"00",
35173=>X"00",
35174=>X"00",
35175=>X"00",
35176=>X"00",
35177=>X"00",
35178=>X"00",
35179=>X"00",
35180=>X"00",
35181=>X"00",
35182=>X"00",
35183=>X"00",
35184=>X"00",
35185=>X"00",
35186=>X"00",
35187=>X"00",
35188=>X"00",
35189=>X"00",
35190=>X"00",
35191=>X"00",
35192=>X"00",
35193=>X"00",
35194=>X"00",
35195=>X"00",
35196=>X"00",
35197=>X"00",
35198=>X"00",
35199=>X"00",
35200=>X"00",
35201=>X"00",
35202=>X"00",
35203=>X"00",
35204=>X"00",
35205=>X"00",
35206=>X"00",
35207=>X"00",
35208=>X"00",
35209=>X"00",
35210=>X"00",
35211=>X"00",
35212=>X"00",
35213=>X"00",
35214=>X"00",
35215=>X"00",
35216=>X"00",
35217=>X"00",
35218=>X"00",
35219=>X"00",
35220=>X"00",
35221=>X"00",
35222=>X"00",
35223=>X"00",
35224=>X"00",
35225=>X"00",
35226=>X"00",
35227=>X"00",
35228=>X"00",
35229=>X"00",
35230=>X"00",
35231=>X"00",
35232=>X"00",
35233=>X"00",
35234=>X"00",
35235=>X"00",
35236=>X"00",
35237=>X"00",
35238=>X"00",
35239=>X"00",
35240=>X"00",
35241=>X"00",
35242=>X"00",
35243=>X"00",
35244=>X"00",
35245=>X"00",
35246=>X"00",
35247=>X"00",
35248=>X"00",
35249=>X"00",
35250=>X"00",
35251=>X"00",
35252=>X"00",
35253=>X"00",
35254=>X"00",
35255=>X"00",
35256=>X"00",
35257=>X"00",
35258=>X"00",
35259=>X"00",
35260=>X"00",
35261=>X"00",
35262=>X"00",
35263=>X"00",
35264=>X"00",
35265=>X"00",
35266=>X"00",
35267=>X"00",
35268=>X"00",
35269=>X"00",
35270=>X"00",
35271=>X"00",
35272=>X"00",
35273=>X"00",
35274=>X"00",
35275=>X"00",
35276=>X"00",
35277=>X"00",
35278=>X"00",
35279=>X"00",
35280=>X"00",
35281=>X"00",
35282=>X"00",
35283=>X"00",
35284=>X"00",
35285=>X"00",
35286=>X"00",
35287=>X"00",
35288=>X"00",
35289=>X"00",
35290=>X"00",
35291=>X"00",
35292=>X"00",
35293=>X"00",
35294=>X"00",
35295=>X"00",
35296=>X"00",
35297=>X"00",
35298=>X"00",
35299=>X"00",
35300=>X"00",
35301=>X"00",
35302=>X"00",
35303=>X"00",
35304=>X"00",
35305=>X"00",
35306=>X"00",
35307=>X"00",
35308=>X"00",
35309=>X"00",
35310=>X"00",
35311=>X"00",
35312=>X"00",
35313=>X"00",
35314=>X"00",
35315=>X"00",
35316=>X"00",
35317=>X"00",
35318=>X"00",
35319=>X"00",
35320=>X"00",
35321=>X"00",
35322=>X"00",
35323=>X"00",
35324=>X"00",
35325=>X"00",
35326=>X"00",
35327=>X"00",
35328=>X"00",
35329=>X"00",
35330=>X"00",
35331=>X"00",
35332=>X"00",
35333=>X"00",
35334=>X"00",
35335=>X"00",
35336=>X"00",
35337=>X"00",
35338=>X"00",
35339=>X"00",
35340=>X"00",
35341=>X"00",
35342=>X"00",
35343=>X"00",
35344=>X"00",
35345=>X"00",
35346=>X"00",
35347=>X"00",
35348=>X"00",
35349=>X"00",
35350=>X"00",
35351=>X"00",
35352=>X"00",
35353=>X"00",
35354=>X"00",
35355=>X"00",
35356=>X"00",
35357=>X"00",
35358=>X"00",
35359=>X"00",
35360=>X"00",
35361=>X"00",
35362=>X"00",
35363=>X"00",
35364=>X"00",
35365=>X"00",
35366=>X"00",
35367=>X"00",
35368=>X"00",
35369=>X"00",
35370=>X"00",
35371=>X"00",
35372=>X"00",
35373=>X"00",
35374=>X"00",
35375=>X"00",
35376=>X"00",
35377=>X"00",
35378=>X"00",
35379=>X"00",
35380=>X"00",
35381=>X"00",
35382=>X"00",
35383=>X"00",
35384=>X"00",
35385=>X"00",
35386=>X"00",
35387=>X"00",
35388=>X"00",
35389=>X"00",
35390=>X"00",
35391=>X"00",
35392=>X"00",
35393=>X"00",
35394=>X"00",
35395=>X"00",
35396=>X"00",
35397=>X"00",
35398=>X"00",
35399=>X"00",
35400=>X"00",
35401=>X"00",
35402=>X"00",
35403=>X"00",
35404=>X"00",
35405=>X"00",
35406=>X"00",
35407=>X"00",
35408=>X"00",
35409=>X"00",
35410=>X"00",
35411=>X"00",
35412=>X"00",
35413=>X"00",
35414=>X"00",
35415=>X"00",
35416=>X"00",
35417=>X"00",
35418=>X"00",
35419=>X"00",
35420=>X"00",
35421=>X"00",
35422=>X"00",
35423=>X"00",
35424=>X"00",
35425=>X"00",
35426=>X"00",
35427=>X"00",
35428=>X"00",
35429=>X"00",
35430=>X"00",
35431=>X"00",
35432=>X"00",
35433=>X"00",
35434=>X"00",
35435=>X"00",
35436=>X"00",
35437=>X"00",
35438=>X"00",
35439=>X"00",
35440=>X"00",
35441=>X"00",
35442=>X"00",
35443=>X"00",
35444=>X"00",
35445=>X"00",
35446=>X"00",
35447=>X"00",
35448=>X"00",
35449=>X"00",
35450=>X"00",
35451=>X"00",
35452=>X"00",
35453=>X"00",
35454=>X"00",
35455=>X"00",
35456=>X"00",
35457=>X"00",
35458=>X"00",
35459=>X"00",
35460=>X"00",
35461=>X"00",
35462=>X"00",
35463=>X"00",
35464=>X"00",
35465=>X"00",
35466=>X"00",
35467=>X"00",
35468=>X"00",
35469=>X"00",
35470=>X"00",
35471=>X"00",
35472=>X"00",
35473=>X"00",
35474=>X"00",
35475=>X"00",
35476=>X"00",
35477=>X"00",
35478=>X"00",
35479=>X"00",
35480=>X"00",
35481=>X"00",
35482=>X"00",
35483=>X"00",
35484=>X"00",
35485=>X"00",
35486=>X"00",
35487=>X"00",
35488=>X"00",
35489=>X"00",
35490=>X"00",
35491=>X"00",
35492=>X"00",
35493=>X"00",
35494=>X"00",
35495=>X"00",
35496=>X"00",
35497=>X"00",
35498=>X"00",
35499=>X"00",
35500=>X"00",
35501=>X"00",
35502=>X"00",
35503=>X"00",
35504=>X"00",
35505=>X"00",
35506=>X"00",
35507=>X"00",
35508=>X"00",
35509=>X"00",
35510=>X"00",
35511=>X"00",
35512=>X"00",
35513=>X"00",
35514=>X"00",
35515=>X"00",
35516=>X"00",
35517=>X"00",
35518=>X"00",
35519=>X"00",
35520=>X"00",
35521=>X"00",
35522=>X"00",
35523=>X"00",
35524=>X"00",
35525=>X"00",
35526=>X"00",
35527=>X"00",
35528=>X"00",
35529=>X"00",
35530=>X"00",
35531=>X"00",
35532=>X"00",
35533=>X"00",
35534=>X"00",
35535=>X"00",
35536=>X"00",
35537=>X"00",
35538=>X"00",
35539=>X"00",
35540=>X"00",
35541=>X"00",
35542=>X"00",
35543=>X"00",
35544=>X"00",
35545=>X"00",
35546=>X"00",
35547=>X"00",
35548=>X"00",
35549=>X"00",
35550=>X"00",
35551=>X"00",
35552=>X"00",
35553=>X"00",
35554=>X"00",
35555=>X"00",
35556=>X"00",
35557=>X"00",
35558=>X"00",
35559=>X"00",
35560=>X"00",
35561=>X"00",
35562=>X"00",
35563=>X"00",
35564=>X"00",
35565=>X"00",
35566=>X"00",
35567=>X"00",
35568=>X"00",
35569=>X"00",
35570=>X"00",
35571=>X"00",
35572=>X"00",
35573=>X"00",
35574=>X"00",
35575=>X"00",
35576=>X"00",
35577=>X"00",
35578=>X"00",
35579=>X"00",
35580=>X"00",
35581=>X"00",
35582=>X"00",
35583=>X"00",
35584=>X"00",
35585=>X"00",
35586=>X"00",
35587=>X"00",
35588=>X"00",
35589=>X"00",
35590=>X"00",
35591=>X"00",
35592=>X"00",
35593=>X"00",
35594=>X"00",
35595=>X"00",
35596=>X"00",
35597=>X"00",
35598=>X"00",
35599=>X"00",
35600=>X"00",
35601=>X"00",
35602=>X"00",
35603=>X"00",
35604=>X"00",
35605=>X"00",
35606=>X"00",
35607=>X"00",
35608=>X"00",
35609=>X"00",
35610=>X"00",
35611=>X"00",
35612=>X"00",
35613=>X"00",
35614=>X"00",
35615=>X"00",
35616=>X"00",
35617=>X"00",
35618=>X"00",
35619=>X"00",
35620=>X"00",
35621=>X"00",
35622=>X"00",
35623=>X"00",
35624=>X"00",
35625=>X"00",
35626=>X"00",
35627=>X"00",
35628=>X"00",
35629=>X"00",
35630=>X"00",
35631=>X"00",
35632=>X"00",
35633=>X"00",
35634=>X"00",
35635=>X"00",
35636=>X"00",
35637=>X"00",
35638=>X"00",
35639=>X"00",
35640=>X"00",
35641=>X"00",
35642=>X"00",
35643=>X"00",
35644=>X"00",
35645=>X"00",
35646=>X"00",
35647=>X"00",
35648=>X"00",
35649=>X"00",
35650=>X"00",
35651=>X"00",
35652=>X"00",
35653=>X"00",
35654=>X"00",
35655=>X"00",
35656=>X"00",
35657=>X"00",
35658=>X"00",
35659=>X"00",
35660=>X"00",
35661=>X"00",
35662=>X"00",
35663=>X"00",
35664=>X"00",
35665=>X"00",
35666=>X"00",
35667=>X"00",
35668=>X"00",
35669=>X"00",
35670=>X"00",
35671=>X"00",
35672=>X"00",
35673=>X"00",
35674=>X"00",
35675=>X"00",
35676=>X"00",
35677=>X"00",
35678=>X"00",
35679=>X"00",
35680=>X"00",
35681=>X"00",
35682=>X"00",
35683=>X"00",
35684=>X"00",
35685=>X"00",
35686=>X"00",
35687=>X"00",
35688=>X"00",
35689=>X"00",
35690=>X"00",
35691=>X"00",
35692=>X"00",
35693=>X"00",
35694=>X"00",
35695=>X"00",
35696=>X"00",
35697=>X"00",
35698=>X"00",
35699=>X"00",
35700=>X"00",
35701=>X"00",
35702=>X"00",
35703=>X"00",
35704=>X"00",
35705=>X"00",
35706=>X"00",
35707=>X"00",
35708=>X"00",
35709=>X"00",
35710=>X"00",
35711=>X"00",
35712=>X"00",
35713=>X"00",
35714=>X"00",
35715=>X"00",
35716=>X"00",
35717=>X"00",
35718=>X"00",
35719=>X"00",
35720=>X"00",
35721=>X"00",
35722=>X"00",
35723=>X"00",
35724=>X"00",
35725=>X"00",
35726=>X"00",
35727=>X"00",
35728=>X"00",
35729=>X"00",
35730=>X"00",
35731=>X"00",
35732=>X"00",
35733=>X"00",
35734=>X"00",
35735=>X"00",
35736=>X"00",
35737=>X"00",
35738=>X"00",
35739=>X"00",
35740=>X"00",
35741=>X"00",
35742=>X"00",
35743=>X"00",
35744=>X"00",
35745=>X"00",
35746=>X"00",
35747=>X"00",
35748=>X"00",
35749=>X"00",
35750=>X"00",
35751=>X"00",
35752=>X"00",
35753=>X"00",
35754=>X"00",
35755=>X"00",
35756=>X"00",
35757=>X"00",
35758=>X"00",
35759=>X"00",
35760=>X"00",
35761=>X"00",
35762=>X"00",
35763=>X"00",
35764=>X"00",
35765=>X"00",
35766=>X"00",
35767=>X"00",
35768=>X"00",
35769=>X"00",
35770=>X"00",
35771=>X"00",
35772=>X"00",
35773=>X"00",
35774=>X"00",
35775=>X"00",
35776=>X"00",
35777=>X"00",
35778=>X"00",
35779=>X"00",
35780=>X"00",
35781=>X"00",
35782=>X"00",
35783=>X"00",
35784=>X"00",
35785=>X"00",
35786=>X"00",
35787=>X"00",
35788=>X"00",
35789=>X"00",
35790=>X"00",
35791=>X"00",
35792=>X"00",
35793=>X"00",
35794=>X"00",
35795=>X"00",
35796=>X"00",
35797=>X"00",
35798=>X"00",
35799=>X"00",
35800=>X"00",
35801=>X"00",
35802=>X"00",
35803=>X"00",
35804=>X"00",
35805=>X"00",
35806=>X"00",
35807=>X"00",
35808=>X"00",
35809=>X"00",
35810=>X"00",
35811=>X"00",
35812=>X"00",
35813=>X"00",
35814=>X"00",
35815=>X"00",
35816=>X"00",
35817=>X"00",
35818=>X"00",
35819=>X"00",
35820=>X"00",
35821=>X"00",
35822=>X"00",
35823=>X"00",
35824=>X"00",
35825=>X"00",
35826=>X"00",
35827=>X"00",
35828=>X"00",
35829=>X"00",
35830=>X"00",
35831=>X"00",
35832=>X"00",
35833=>X"00",
35834=>X"00",
35835=>X"00",
35836=>X"00",
35837=>X"00",
35838=>X"00",
35839=>X"00",
35840=>X"00",
35841=>X"00",
35842=>X"00",
35843=>X"00",
35844=>X"00",
35845=>X"00",
35846=>X"00",
35847=>X"00",
35848=>X"00",
35849=>X"00",
35850=>X"00",
35851=>X"00",
35852=>X"00",
35853=>X"00",
35854=>X"00",
35855=>X"00",
35856=>X"00",
35857=>X"00",
35858=>X"00",
35859=>X"00",
35860=>X"00",
35861=>X"00",
35862=>X"00",
35863=>X"00",
35864=>X"00",
35865=>X"00",
35866=>X"00",
35867=>X"00",
35868=>X"00",
35869=>X"00",
35870=>X"00",
35871=>X"00",
35872=>X"00",
35873=>X"00",
35874=>X"00",
35875=>X"00",
35876=>X"00",
35877=>X"00",
35878=>X"00",
35879=>X"00",
35880=>X"00",
35881=>X"00",
35882=>X"00",
35883=>X"00",
35884=>X"00",
35885=>X"00",
35886=>X"00",
35887=>X"00",
35888=>X"00",
35889=>X"00",
35890=>X"00",
35891=>X"00",
35892=>X"00",
35893=>X"00",
35894=>X"00",
35895=>X"00",
35896=>X"00",
35897=>X"00",
35898=>X"00",
35899=>X"00",
35900=>X"00",
35901=>X"00",
35902=>X"00",
35903=>X"00",
35904=>X"00",
35905=>X"00",
35906=>X"00",
35907=>X"00",
35908=>X"00",
35909=>X"00",
35910=>X"00",
35911=>X"00",
35912=>X"00",
35913=>X"00",
35914=>X"00",
35915=>X"00",
35916=>X"00",
35917=>X"00",
35918=>X"00",
35919=>X"00",
35920=>X"00",
35921=>X"00",
35922=>X"00",
35923=>X"00",
35924=>X"00",
35925=>X"00",
35926=>X"00",
35927=>X"00",
35928=>X"00",
35929=>X"00",
35930=>X"00",
35931=>X"00",
35932=>X"00",
35933=>X"00",
35934=>X"00",
35935=>X"00",
35936=>X"00",
35937=>X"00",
35938=>X"00",
35939=>X"00",
35940=>X"00",
35941=>X"00",
35942=>X"00",
35943=>X"00",
35944=>X"00",
35945=>X"00",
35946=>X"00",
35947=>X"00",
35948=>X"00",
35949=>X"00",
35950=>X"00",
35951=>X"00",
35952=>X"00",
35953=>X"00",
35954=>X"00",
35955=>X"00",
35956=>X"00",
35957=>X"00",
35958=>X"00",
35959=>X"00",
35960=>X"00",
35961=>X"00",
35962=>X"00",
35963=>X"00",
35964=>X"00",
35965=>X"00",
35966=>X"00",
35967=>X"00",
35968=>X"00",
35969=>X"00",
35970=>X"00",
35971=>X"00",
35972=>X"00",
35973=>X"00",
35974=>X"00",
35975=>X"00",
35976=>X"00",
35977=>X"00",
35978=>X"00",
35979=>X"00",
35980=>X"00",
35981=>X"00",
35982=>X"00",
35983=>X"00",
35984=>X"00",
35985=>X"00",
35986=>X"00",
35987=>X"00",
35988=>X"00",
35989=>X"00",
35990=>X"00",
35991=>X"00",
35992=>X"00",
35993=>X"00",
35994=>X"00",
35995=>X"00",
35996=>X"00",
35997=>X"00",
35998=>X"00",
35999=>X"00",
36000=>X"00",
36001=>X"00",
36002=>X"00",
36003=>X"00",
36004=>X"00",
36005=>X"00",
36006=>X"00",
36007=>X"00",
36008=>X"00",
36009=>X"00",
36010=>X"00",
36011=>X"00",
36012=>X"00",
36013=>X"00",
36014=>X"00",
36015=>X"00",
36016=>X"00",
36017=>X"00",
36018=>X"00",
36019=>X"00",
36020=>X"00",
36021=>X"00",
36022=>X"00",
36023=>X"00",
36024=>X"00",
36025=>X"00",
36026=>X"00",
36027=>X"00",
36028=>X"00",
36029=>X"00",
36030=>X"00",
36031=>X"00",
36032=>X"00",
36033=>X"00",
36034=>X"00",
36035=>X"00",
36036=>X"00",
36037=>X"00",
36038=>X"00",
36039=>X"00",
36040=>X"00",
36041=>X"00",
36042=>X"00",
36043=>X"00",
36044=>X"00",
36045=>X"00",
36046=>X"00",
36047=>X"00",
36048=>X"00",
36049=>X"00",
36050=>X"00",
36051=>X"00",
36052=>X"00",
36053=>X"00",
36054=>X"00",
36055=>X"00",
36056=>X"00",
36057=>X"00",
36058=>X"00",
36059=>X"00",
36060=>X"00",
36061=>X"00",
36062=>X"00",
36063=>X"00",
36064=>X"00",
36065=>X"00",
36066=>X"00",
36067=>X"00",
36068=>X"00",
36069=>X"00",
36070=>X"00",
36071=>X"00",
36072=>X"00",
36073=>X"00",
36074=>X"00",
36075=>X"00",
36076=>X"00",
36077=>X"00",
36078=>X"00",
36079=>X"00",
36080=>X"00",
36081=>X"00",
36082=>X"00",
36083=>X"00",
36084=>X"00",
36085=>X"00",
36086=>X"00",
36087=>X"00",
36088=>X"00",
36089=>X"00",
36090=>X"00",
36091=>X"00",
36092=>X"00",
36093=>X"00",
36094=>X"00",
36095=>X"00",
36096=>X"00",
36097=>X"00",
36098=>X"00",
36099=>X"00",
36100=>X"00",
36101=>X"00",
36102=>X"00",
36103=>X"00",
36104=>X"00",
36105=>X"00",
36106=>X"00",
36107=>X"00",
36108=>X"00",
36109=>X"00",
36110=>X"00",
36111=>X"00",
36112=>X"00",
36113=>X"00",
36114=>X"00",
36115=>X"00",
36116=>X"00",
36117=>X"00",
36118=>X"00",
36119=>X"00",
36120=>X"00",
36121=>X"00",
36122=>X"00",
36123=>X"00",
36124=>X"00",
36125=>X"00",
36126=>X"00",
36127=>X"00",
36128=>X"00",
36129=>X"00",
36130=>X"00",
36131=>X"00",
36132=>X"00",
36133=>X"00",
36134=>X"00",
36135=>X"00",
36136=>X"00",
36137=>X"00",
36138=>X"00",
36139=>X"00",
36140=>X"00",
36141=>X"00",
36142=>X"00",
36143=>X"00",
36144=>X"00",
36145=>X"00",
36146=>X"00",
36147=>X"00",
36148=>X"00",
36149=>X"00",
36150=>X"00",
36151=>X"00",
36152=>X"00",
36153=>X"00",
36154=>X"00",
36155=>X"00",
36156=>X"00",
36157=>X"00",
36158=>X"00",
36159=>X"00",
36160=>X"00",
36161=>X"00",
36162=>X"00",
36163=>X"00",
36164=>X"00",
36165=>X"00",
36166=>X"00",
36167=>X"00",
36168=>X"00",
36169=>X"00",
36170=>X"00",
36171=>X"00",
36172=>X"00",
36173=>X"00",
36174=>X"00",
36175=>X"00",
36176=>X"00",
36177=>X"00",
36178=>X"00",
36179=>X"00",
36180=>X"00",
36181=>X"00",
36182=>X"00",
36183=>X"00",
36184=>X"00",
36185=>X"00",
36186=>X"00",
36187=>X"00",
36188=>X"00",
36189=>X"00",
36190=>X"00",
36191=>X"00",
36192=>X"00",
36193=>X"00",
36194=>X"00",
36195=>X"00",
36196=>X"00",
36197=>X"00",
36198=>X"00",
36199=>X"00",
36200=>X"00",
36201=>X"00",
36202=>X"00",
36203=>X"00",
36204=>X"00",
36205=>X"00",
36206=>X"00",
36207=>X"00",
36208=>X"00",
36209=>X"00",
36210=>X"00",
36211=>X"00",
36212=>X"00",
36213=>X"00",
36214=>X"00",
36215=>X"00",
36216=>X"00",
36217=>X"00",
36218=>X"00",
36219=>X"00",
36220=>X"00",
36221=>X"00",
36222=>X"00",
36223=>X"00",
36224=>X"00",
36225=>X"00",
36226=>X"00",
36227=>X"00",
36228=>X"00",
36229=>X"00",
36230=>X"00",
36231=>X"00",
36232=>X"00",
36233=>X"00",
36234=>X"00",
36235=>X"00",
36236=>X"00",
36237=>X"00",
36238=>X"00",
36239=>X"00",
36240=>X"00",
36241=>X"00",
36242=>X"00",
36243=>X"00",
36244=>X"00",
36245=>X"00",
36246=>X"00",
36247=>X"00",
36248=>X"00",
36249=>X"00",
36250=>X"00",
36251=>X"00",
36252=>X"00",
36253=>X"00",
36254=>X"00",
36255=>X"00",
36256=>X"00",
36257=>X"00",
36258=>X"00",
36259=>X"00",
36260=>X"00",
36261=>X"00",
36262=>X"00",
36263=>X"00",
36264=>X"00",
36265=>X"00",
36266=>X"00",
36267=>X"00",
36268=>X"00",
36269=>X"00",
36270=>X"00",
36271=>X"00",
36272=>X"00",
36273=>X"00",
36274=>X"00",
36275=>X"00",
36276=>X"00",
36277=>X"00",
36278=>X"00",
36279=>X"00",
36280=>X"00",
36281=>X"00",
36282=>X"00",
36283=>X"00",
36284=>X"00",
36285=>X"00",
36286=>X"00",
36287=>X"00",
36288=>X"00",
36289=>X"00",
36290=>X"00",
36291=>X"00",
36292=>X"00",
36293=>X"00",
36294=>X"00",
36295=>X"00",
36296=>X"00",
36297=>X"00",
36298=>X"00",
36299=>X"00",
36300=>X"00",
36301=>X"00",
36302=>X"00",
36303=>X"00",
36304=>X"00",
36305=>X"00",
36306=>X"00",
36307=>X"00",
36308=>X"00",
36309=>X"00",
36310=>X"00",
36311=>X"00",
36312=>X"00",
36313=>X"00",
36314=>X"00",
36315=>X"00",
36316=>X"00",
36317=>X"00",
36318=>X"00",
36319=>X"00",
36320=>X"00",
36321=>X"00",
36322=>X"00",
36323=>X"00",
36324=>X"00",
36325=>X"00",
36326=>X"00",
36327=>X"00",
36328=>X"00",
36329=>X"00",
36330=>X"00",
36331=>X"00",
36332=>X"00",
36333=>X"00",
36334=>X"00",
36335=>X"00",
36336=>X"00",
36337=>X"00",
36338=>X"00",
36339=>X"00",
36340=>X"00",
36341=>X"00",
36342=>X"00",
36343=>X"00",
36344=>X"00",
36345=>X"00",
36346=>X"00",
36347=>X"00",
36348=>X"00",
36349=>X"00",
36350=>X"00",
36351=>X"00",
36352=>X"00",
36353=>X"00",
36354=>X"00",
36355=>X"00",
36356=>X"00",
36357=>X"00",
36358=>X"00",
36359=>X"00",
36360=>X"00",
36361=>X"00",
36362=>X"00",
36363=>X"00",
36364=>X"00",
36365=>X"00",
36366=>X"00",
36367=>X"00",
36368=>X"00",
36369=>X"00",
36370=>X"00",
36371=>X"00",
36372=>X"00",
36373=>X"00",
36374=>X"00",
36375=>X"00",
36376=>X"00",
36377=>X"00",
36378=>X"00",
36379=>X"00",
36380=>X"00",
36381=>X"00",
36382=>X"00",
36383=>X"00",
36384=>X"00",
36385=>X"00",
36386=>X"00",
36387=>X"00",
36388=>X"00",
36389=>X"00",
36390=>X"00",
36391=>X"00",
36392=>X"00",
36393=>X"00",
36394=>X"00",
36395=>X"00",
36396=>X"00",
36397=>X"00",
36398=>X"00",
36399=>X"00",
36400=>X"00",
36401=>X"00",
36402=>X"00",
36403=>X"00",
36404=>X"00",
36405=>X"00",
36406=>X"00",
36407=>X"00",
36408=>X"00",
36409=>X"00",
36410=>X"00",
36411=>X"00",
36412=>X"00",
36413=>X"00",
36414=>X"00",
36415=>X"00",
36416=>X"00",
36417=>X"00",
36418=>X"00",
36419=>X"00",
36420=>X"00",
36421=>X"00",
36422=>X"00",
36423=>X"00",
36424=>X"00",
36425=>X"00",
36426=>X"00",
36427=>X"00",
36428=>X"00",
36429=>X"00",
36430=>X"00",
36431=>X"00",
36432=>X"00",
36433=>X"00",
36434=>X"00",
36435=>X"00",
36436=>X"00",
36437=>X"00",
36438=>X"00",
36439=>X"00",
36440=>X"00",
36441=>X"00",
36442=>X"00",
36443=>X"00",
36444=>X"00",
36445=>X"00",
36446=>X"00",
36447=>X"00",
36448=>X"00",
36449=>X"00",
36450=>X"00",
36451=>X"00",
36452=>X"00",
36453=>X"00",
36454=>X"00",
36455=>X"00",
36456=>X"00",
36457=>X"00",
36458=>X"00",
36459=>X"00",
36460=>X"00",
36461=>X"00",
36462=>X"00",
36463=>X"00",
36464=>X"00",
36465=>X"00",
36466=>X"00",
36467=>X"00",
36468=>X"00",
36469=>X"00",
36470=>X"00",
36471=>X"00",
36472=>X"00",
36473=>X"00",
36474=>X"00",
36475=>X"00",
36476=>X"00",
36477=>X"00",
36478=>X"00",
36479=>X"00",
36480=>X"00",
36481=>X"00",
36482=>X"00",
36483=>X"00",
36484=>X"00",
36485=>X"00",
36486=>X"00",
36487=>X"00",
36488=>X"00",
36489=>X"00",
36490=>X"00",
36491=>X"00",
36492=>X"00",
36493=>X"00",
36494=>X"00",
36495=>X"00",
36496=>X"00",
36497=>X"00",
36498=>X"00",
36499=>X"00",
36500=>X"00",
36501=>X"00",
36502=>X"00",
36503=>X"00",
36504=>X"00",
36505=>X"00",
36506=>X"00",
36507=>X"00",
36508=>X"00",
36509=>X"00",
36510=>X"00",
36511=>X"00",
36512=>X"00",
36513=>X"00",
36514=>X"00",
36515=>X"00",
36516=>X"00",
36517=>X"00",
36518=>X"00",
36519=>X"00",
36520=>X"00",
36521=>X"00",
36522=>X"00",
36523=>X"00",
36524=>X"00",
36525=>X"00",
36526=>X"00",
36527=>X"00",
36528=>X"00",
36529=>X"00",
36530=>X"00",
36531=>X"00",
36532=>X"00",
36533=>X"00",
36534=>X"00",
36535=>X"00",
36536=>X"00",
36537=>X"00",
36538=>X"00",
36539=>X"00",
36540=>X"00",
36541=>X"00",
36542=>X"00",
36543=>X"00",
36544=>X"00",
36545=>X"00",
36546=>X"00",
36547=>X"00",
36548=>X"00",
36549=>X"00",
36550=>X"00",
36551=>X"00",
36552=>X"00",
36553=>X"00",
36554=>X"00",
36555=>X"00",
36556=>X"00",
36557=>X"00",
36558=>X"00",
36559=>X"00",
36560=>X"00",
36561=>X"00",
36562=>X"00",
36563=>X"00",
36564=>X"00",
36565=>X"00",
36566=>X"00",
36567=>X"00",
36568=>X"00",
36569=>X"00",
36570=>X"00",
36571=>X"00",
36572=>X"00",
36573=>X"00",
36574=>X"00",
36575=>X"00",
36576=>X"00",
36577=>X"00",
36578=>X"00",
36579=>X"00",
36580=>X"00",
36581=>X"00",
36582=>X"00",
36583=>X"00",
36584=>X"00",
36585=>X"00",
36586=>X"00",
36587=>X"00",
36588=>X"00",
36589=>X"00",
36590=>X"00",
36591=>X"00",
36592=>X"00",
36593=>X"00",
36594=>X"00",
36595=>X"00",
36596=>X"00",
36597=>X"00",
36598=>X"00",
36599=>X"00",
36600=>X"00",
36601=>X"00",
36602=>X"00",
36603=>X"00",
36604=>X"00",
36605=>X"00",
36606=>X"00",
36607=>X"00",
36608=>X"00",
36609=>X"00",
36610=>X"00",
36611=>X"00",
36612=>X"00",
36613=>X"00",
36614=>X"00",
36615=>X"00",
36616=>X"00",
36617=>X"00",
36618=>X"00",
36619=>X"00",
36620=>X"00",
36621=>X"00",
36622=>X"00",
36623=>X"00",
36624=>X"00",
36625=>X"00",
36626=>X"00",
36627=>X"00",
36628=>X"00",
36629=>X"00",
36630=>X"00",
36631=>X"00",
36632=>X"00",
36633=>X"00",
36634=>X"00",
36635=>X"00",
36636=>X"00",
36637=>X"00",
36638=>X"00",
36639=>X"00",
36640=>X"00",
36641=>X"00",
36642=>X"00",
36643=>X"00",
36644=>X"00",
36645=>X"00",
36646=>X"00",
36647=>X"00",
36648=>X"00",
36649=>X"00",
36650=>X"00",
36651=>X"00",
36652=>X"00",
36653=>X"00",
36654=>X"00",
36655=>X"00",
36656=>X"00",
36657=>X"00",
36658=>X"00",
36659=>X"00",
36660=>X"00",
36661=>X"00",
36662=>X"00",
36663=>X"00",
36664=>X"00",
36665=>X"00",
36666=>X"00",
36667=>X"00",
36668=>X"00",
36669=>X"00",
36670=>X"00",
36671=>X"00",
36672=>X"00",
36673=>X"00",
36674=>X"00",
36675=>X"00",
36676=>X"00",
36677=>X"00",
36678=>X"00",
36679=>X"00",
36680=>X"00",
36681=>X"00",
36682=>X"00",
36683=>X"00",
36684=>X"00",
36685=>X"00",
36686=>X"00",
36687=>X"00",
36688=>X"00",
36689=>X"00",
36690=>X"00",
36691=>X"00",
36692=>X"00",
36693=>X"00",
36694=>X"00",
36695=>X"00",
36696=>X"00",
36697=>X"00",
36698=>X"00",
36699=>X"00",
36700=>X"00",
36701=>X"00",
36702=>X"00",
36703=>X"00",
36704=>X"00",
36705=>X"00",
36706=>X"00",
36707=>X"00",
36708=>X"00",
36709=>X"00",
36710=>X"00",
36711=>X"00",
36712=>X"00",
36713=>X"00",
36714=>X"00",
36715=>X"00",
36716=>X"00",
36717=>X"00",
36718=>X"00",
36719=>X"00",
36720=>X"00",
36721=>X"00",
36722=>X"00",
36723=>X"00",
36724=>X"00",
36725=>X"00",
36726=>X"00",
36727=>X"00",
36728=>X"00",
36729=>X"00",
36730=>X"00",
36731=>X"00",
36732=>X"00",
36733=>X"00",
36734=>X"00",
36735=>X"00",
36736=>X"00",
36737=>X"00",
36738=>X"00",
36739=>X"00",
36740=>X"00",
36741=>X"00",
36742=>X"00",
36743=>X"00",
36744=>X"00",
36745=>X"00",
36746=>X"00",
36747=>X"00",
36748=>X"00",
36749=>X"00",
36750=>X"00",
36751=>X"00",
36752=>X"00",
36753=>X"00",
36754=>X"00",
36755=>X"00",
36756=>X"00",
36757=>X"00",
36758=>X"00",
36759=>X"00",
36760=>X"00",
36761=>X"00",
36762=>X"00",
36763=>X"00",
36764=>X"00",
36765=>X"00",
36766=>X"00",
36767=>X"00",
36768=>X"00",
36769=>X"00",
36770=>X"00",
36771=>X"00",
36772=>X"00",
36773=>X"00",
36774=>X"00",
36775=>X"00",
36776=>X"00",
36777=>X"00",
36778=>X"00",
36779=>X"00",
36780=>X"00",
36781=>X"00",
36782=>X"00",
36783=>X"00",
36784=>X"00",
36785=>X"00",
36786=>X"00",
36787=>X"00",
36788=>X"00",
36789=>X"00",
36790=>X"00",
36791=>X"00",
36792=>X"00",
36793=>X"00",
36794=>X"00",
36795=>X"00",
36796=>X"00",
36797=>X"00",
36798=>X"00",
36799=>X"00",
36800=>X"00",
36801=>X"00",
36802=>X"00",
36803=>X"00",
36804=>X"00",
36805=>X"00",
36806=>X"00",
36807=>X"00",
36808=>X"00",
36809=>X"00",
36810=>X"00",
36811=>X"00",
36812=>X"00",
36813=>X"00",
36814=>X"00",
36815=>X"00",
36816=>X"00",
36817=>X"00",
36818=>X"00",
36819=>X"00",
36820=>X"00",
36821=>X"00",
36822=>X"00",
36823=>X"00",
36824=>X"00",
36825=>X"00",
36826=>X"00",
36827=>X"00",
36828=>X"00",
36829=>X"00",
36830=>X"00",
36831=>X"00",
36832=>X"00",
36833=>X"00",
36834=>X"00",
36835=>X"00",
36836=>X"00",
36837=>X"00",
36838=>X"00",
36839=>X"00",
36840=>X"00",
36841=>X"00",
36842=>X"00",
36843=>X"00",
36844=>X"00",
36845=>X"00",
36846=>X"00",
36847=>X"00",
36848=>X"00",
36849=>X"00",
36850=>X"00",
36851=>X"00",
36852=>X"00",
36853=>X"00",
36854=>X"00",
36855=>X"00",
36856=>X"00",
36857=>X"00",
36858=>X"00",
36859=>X"00",
36860=>X"00",
36861=>X"00",
36862=>X"00",
36863=>X"00",
36864=>X"00",
36865=>X"00",
36866=>X"00",
36867=>X"00",
36868=>X"00",
36869=>X"00",
36870=>X"00",
36871=>X"00",
36872=>X"00",
36873=>X"00",
36874=>X"00",
36875=>X"00",
36876=>X"00",
36877=>X"00",
36878=>X"00",
36879=>X"00",
36880=>X"00",
36881=>X"00",
36882=>X"00",
36883=>X"00",
36884=>X"00",
36885=>X"00",
36886=>X"00",
36887=>X"00",
36888=>X"00",
36889=>X"00",
36890=>X"00",
36891=>X"00",
36892=>X"00",
36893=>X"00",
36894=>X"00",
36895=>X"00",
36896=>X"00",
36897=>X"00",
36898=>X"00",
36899=>X"00",
36900=>X"00",
36901=>X"00",
36902=>X"00",
36903=>X"00",
36904=>X"00",
36905=>X"00",
36906=>X"00",
36907=>X"00",
36908=>X"00",
36909=>X"00",
36910=>X"00",
36911=>X"00",
36912=>X"00",
36913=>X"00",
36914=>X"00",
36915=>X"00",
36916=>X"00",
36917=>X"00",
36918=>X"00",
36919=>X"00",
36920=>X"00",
36921=>X"00",
36922=>X"00",
36923=>X"00",
36924=>X"00",
36925=>X"00",
36926=>X"00",
36927=>X"00",
36928=>X"00",
36929=>X"00",
36930=>X"00",
36931=>X"00",
36932=>X"00",
36933=>X"00",
36934=>X"00",
36935=>X"00",
36936=>X"00",
36937=>X"00",
36938=>X"00",
36939=>X"00",
36940=>X"00",
36941=>X"00",
36942=>X"00",
36943=>X"00",
36944=>X"00",
36945=>X"00",
36946=>X"00",
36947=>X"00",
36948=>X"00",
36949=>X"00",
36950=>X"00",
36951=>X"00",
36952=>X"00",
36953=>X"00",
36954=>X"00",
36955=>X"00",
36956=>X"00",
36957=>X"00",
36958=>X"00",
36959=>X"00",
36960=>X"00",
36961=>X"00",
36962=>X"00",
36963=>X"00",
36964=>X"00",
36965=>X"00",
36966=>X"00",
36967=>X"00",
36968=>X"00",
36969=>X"00",
36970=>X"00",
36971=>X"00",
36972=>X"00",
36973=>X"00",
36974=>X"00",
36975=>X"00",
36976=>X"00",
36977=>X"00",
36978=>X"00",
36979=>X"00",
36980=>X"00",
36981=>X"00",
36982=>X"00",
36983=>X"00",
36984=>X"00",
36985=>X"00",
36986=>X"00",
36987=>X"00",
36988=>X"00",
36989=>X"00",
36990=>X"00",
36991=>X"00",
36992=>X"00",
36993=>X"00",
36994=>X"00",
36995=>X"00",
36996=>X"00",
36997=>X"00",
36998=>X"00",
36999=>X"00",
37000=>X"00",
37001=>X"00",
37002=>X"00",
37003=>X"00",
37004=>X"00",
37005=>X"00",
37006=>X"00",
37007=>X"00",
37008=>X"00",
37009=>X"00",
37010=>X"00",
37011=>X"00",
37012=>X"00",
37013=>X"00",
37014=>X"00",
37015=>X"00",
37016=>X"00",
37017=>X"00",
37018=>X"00",
37019=>X"00",
37020=>X"00",
37021=>X"00",
37022=>X"00",
37023=>X"00",
37024=>X"00",
37025=>X"00",
37026=>X"00",
37027=>X"00",
37028=>X"00",
37029=>X"00",
37030=>X"00",
37031=>X"00",
37032=>X"00",
37033=>X"00",
37034=>X"00",
37035=>X"00",
37036=>X"00",
37037=>X"00",
37038=>X"00",
37039=>X"00",
37040=>X"00",
37041=>X"00",
37042=>X"00",
37043=>X"00",
37044=>X"00",
37045=>X"00",
37046=>X"00",
37047=>X"00",
37048=>X"00",
37049=>X"00",
37050=>X"00",
37051=>X"00",
37052=>X"00",
37053=>X"00",
37054=>X"00",
37055=>X"00",
37056=>X"00",
37057=>X"00",
37058=>X"00",
37059=>X"00",
37060=>X"00",
37061=>X"00",
37062=>X"00",
37063=>X"00",
37064=>X"00",
37065=>X"00",
37066=>X"00",
37067=>X"00",
37068=>X"00",
37069=>X"00",
37070=>X"00",
37071=>X"00",
37072=>X"00",
37073=>X"00",
37074=>X"00",
37075=>X"00",
37076=>X"00",
37077=>X"00",
37078=>X"00",
37079=>X"00",
37080=>X"00",
37081=>X"00",
37082=>X"00",
37083=>X"00",
37084=>X"00",
37085=>X"00",
37086=>X"00",
37087=>X"00",
37088=>X"00",
37089=>X"00",
37090=>X"00",
37091=>X"00",
37092=>X"00",
37093=>X"00",
37094=>X"00",
37095=>X"00",
37096=>X"00",
37097=>X"00",
37098=>X"00",
37099=>X"00",
37100=>X"00",
37101=>X"00",
37102=>X"00",
37103=>X"00",
37104=>X"00",
37105=>X"00",
37106=>X"00",
37107=>X"00",
37108=>X"00",
37109=>X"00",
37110=>X"00",
37111=>X"00",
37112=>X"00",
37113=>X"00",
37114=>X"00",
37115=>X"00",
37116=>X"00",
37117=>X"00",
37118=>X"00",
37119=>X"00",
37120=>X"00",
37121=>X"00",
37122=>X"00",
37123=>X"00",
37124=>X"00",
37125=>X"00",
37126=>X"00",
37127=>X"00",
37128=>X"00",
37129=>X"00",
37130=>X"00",
37131=>X"00",
37132=>X"00",
37133=>X"00",
37134=>X"00",
37135=>X"00",
37136=>X"00",
37137=>X"00",
37138=>X"00",
37139=>X"00",
37140=>X"00",
37141=>X"00",
37142=>X"00",
37143=>X"00",
37144=>X"00",
37145=>X"00",
37146=>X"00",
37147=>X"00",
37148=>X"00",
37149=>X"00",
37150=>X"00",
37151=>X"00",
37152=>X"00",
37153=>X"00",
37154=>X"00",
37155=>X"00",
37156=>X"00",
37157=>X"00",
37158=>X"00",
37159=>X"00",
37160=>X"00",
37161=>X"00",
37162=>X"00",
37163=>X"00",
37164=>X"00",
37165=>X"00",
37166=>X"00",
37167=>X"00",
37168=>X"00",
37169=>X"00",
37170=>X"00",
37171=>X"00",
37172=>X"00",
37173=>X"00",
37174=>X"00",
37175=>X"00",
37176=>X"00",
37177=>X"00",
37178=>X"00",
37179=>X"00",
37180=>X"00",
37181=>X"00",
37182=>X"00",
37183=>X"00",
37184=>X"00",
37185=>X"00",
37186=>X"00",
37187=>X"00",
37188=>X"00",
37189=>X"00",
37190=>X"00",
37191=>X"00",
37192=>X"00",
37193=>X"00",
37194=>X"00",
37195=>X"00",
37196=>X"00",
37197=>X"00",
37198=>X"00",
37199=>X"00",
37200=>X"00",
37201=>X"00",
37202=>X"00",
37203=>X"00",
37204=>X"00",
37205=>X"00",
37206=>X"00",
37207=>X"00",
37208=>X"00",
37209=>X"00",
37210=>X"00",
37211=>X"00",
37212=>X"00",
37213=>X"00",
37214=>X"00",
37215=>X"00",
37216=>X"00",
37217=>X"00",
37218=>X"00",
37219=>X"00",
37220=>X"00",
37221=>X"00",
37222=>X"00",
37223=>X"00",
37224=>X"00",
37225=>X"00",
37226=>X"00",
37227=>X"00",
37228=>X"00",
37229=>X"00",
37230=>X"00",
37231=>X"00",
37232=>X"00",
37233=>X"00",
37234=>X"00",
37235=>X"00",
37236=>X"00",
37237=>X"00",
37238=>X"00",
37239=>X"00",
37240=>X"00",
37241=>X"00",
37242=>X"00",
37243=>X"00",
37244=>X"00",
37245=>X"00",
37246=>X"00",
37247=>X"00",
37248=>X"00",
37249=>X"00",
37250=>X"00",
37251=>X"00",
37252=>X"00",
37253=>X"00",
37254=>X"00",
37255=>X"00",
37256=>X"00",
37257=>X"00",
37258=>X"00",
37259=>X"00",
37260=>X"00",
37261=>X"00",
37262=>X"00",
37263=>X"00",
37264=>X"00",
37265=>X"00",
37266=>X"00",
37267=>X"00",
37268=>X"00",
37269=>X"00",
37270=>X"00",
37271=>X"00",
37272=>X"00",
37273=>X"00",
37274=>X"00",
37275=>X"00",
37276=>X"00",
37277=>X"00",
37278=>X"00",
37279=>X"00",
37280=>X"00",
37281=>X"00",
37282=>X"00",
37283=>X"00",
37284=>X"00",
37285=>X"00",
37286=>X"00",
37287=>X"00",
37288=>X"00",
37289=>X"00",
37290=>X"00",
37291=>X"00",
37292=>X"00",
37293=>X"00",
37294=>X"00",
37295=>X"00",
37296=>X"00",
37297=>X"00",
37298=>X"00",
37299=>X"00",
37300=>X"00",
37301=>X"00",
37302=>X"00",
37303=>X"00",
37304=>X"00",
37305=>X"00",
37306=>X"00",
37307=>X"00",
37308=>X"00",
37309=>X"00",
37310=>X"00",
37311=>X"00",
37312=>X"00",
37313=>X"00",
37314=>X"00",
37315=>X"00",
37316=>X"00",
37317=>X"00",
37318=>X"00",
37319=>X"00",
37320=>X"00",
37321=>X"00",
37322=>X"00",
37323=>X"00",
37324=>X"00",
37325=>X"00",
37326=>X"00",
37327=>X"00",
37328=>X"00",
37329=>X"00",
37330=>X"00",
37331=>X"00",
37332=>X"00",
37333=>X"00",
37334=>X"00",
37335=>X"00",
37336=>X"00",
37337=>X"00",
37338=>X"00",
37339=>X"00",
37340=>X"00",
37341=>X"00",
37342=>X"00",
37343=>X"00",
37344=>X"00",
37345=>X"00",
37346=>X"00",
37347=>X"00",
37348=>X"00",
37349=>X"00",
37350=>X"00",
37351=>X"00",
37352=>X"00",
37353=>X"00",
37354=>X"00",
37355=>X"00",
37356=>X"00",
37357=>X"00",
37358=>X"00",
37359=>X"00",
37360=>X"00",
37361=>X"00",
37362=>X"00",
37363=>X"00",
37364=>X"00",
37365=>X"00",
37366=>X"00",
37367=>X"00",
37368=>X"00",
37369=>X"00",
37370=>X"00",
37371=>X"00",
37372=>X"00",
37373=>X"00",
37374=>X"00",
37375=>X"00",
37376=>X"00",
37377=>X"00",
37378=>X"00",
37379=>X"00",
37380=>X"00",
37381=>X"00",
37382=>X"00",
37383=>X"00",
37384=>X"00",
37385=>X"00",
37386=>X"00",
37387=>X"00",
37388=>X"00",
37389=>X"00",
37390=>X"00",
37391=>X"00",
37392=>X"00",
37393=>X"00",
37394=>X"00",
37395=>X"00",
37396=>X"00",
37397=>X"00",
37398=>X"00",
37399=>X"00",
37400=>X"00",
37401=>X"00",
37402=>X"00",
37403=>X"00",
37404=>X"00",
37405=>X"00",
37406=>X"00",
37407=>X"00",
37408=>X"00",
37409=>X"00",
37410=>X"00",
37411=>X"00",
37412=>X"00",
37413=>X"00",
37414=>X"00",
37415=>X"00",
37416=>X"00",
37417=>X"00",
37418=>X"00",
37419=>X"00",
37420=>X"00",
37421=>X"00",
37422=>X"00",
37423=>X"00",
37424=>X"00",
37425=>X"00",
37426=>X"00",
37427=>X"00",
37428=>X"00",
37429=>X"00",
37430=>X"00",
37431=>X"00",
37432=>X"00",
37433=>X"00",
37434=>X"00",
37435=>X"00",
37436=>X"00",
37437=>X"00",
37438=>X"00",
37439=>X"00",
37440=>X"00",
37441=>X"00",
37442=>X"00",
37443=>X"00",
37444=>X"00",
37445=>X"00",
37446=>X"00",
37447=>X"00",
37448=>X"00",
37449=>X"00",
37450=>X"00",
37451=>X"00",
37452=>X"00",
37453=>X"00",
37454=>X"00",
37455=>X"00",
37456=>X"00",
37457=>X"00",
37458=>X"00",
37459=>X"00",
37460=>X"00",
37461=>X"00",
37462=>X"00",
37463=>X"00",
37464=>X"00",
37465=>X"00",
37466=>X"00",
37467=>X"00",
37468=>X"00",
37469=>X"00",
37470=>X"00",
37471=>X"00",
37472=>X"00",
37473=>X"00",
37474=>X"00",
37475=>X"00",
37476=>X"00",
37477=>X"00",
37478=>X"00",
37479=>X"00",
37480=>X"00",
37481=>X"00",
37482=>X"00",
37483=>X"00",
37484=>X"00",
37485=>X"00",
37486=>X"00",
37487=>X"00",
37488=>X"00",
37489=>X"00",
37490=>X"00",
37491=>X"00",
37492=>X"00",
37493=>X"00",
37494=>X"00",
37495=>X"00",
37496=>X"00",
37497=>X"00",
37498=>X"00",
37499=>X"00",
37500=>X"00",
37501=>X"00",
37502=>X"00",
37503=>X"00",
37504=>X"00",
37505=>X"00",
37506=>X"00",
37507=>X"00",
37508=>X"00",
37509=>X"00",
37510=>X"00",
37511=>X"00",
37512=>X"00",
37513=>X"00",
37514=>X"00",
37515=>X"00",
37516=>X"00",
37517=>X"00",
37518=>X"00",
37519=>X"00",
37520=>X"00",
37521=>X"00",
37522=>X"00",
37523=>X"00",
37524=>X"00",
37525=>X"00",
37526=>X"00",
37527=>X"00",
37528=>X"00",
37529=>X"00",
37530=>X"00",
37531=>X"00",
37532=>X"00",
37533=>X"00",
37534=>X"00",
37535=>X"00",
37536=>X"00",
37537=>X"00",
37538=>X"00",
37539=>X"00",
37540=>X"00",
37541=>X"00",
37542=>X"00",
37543=>X"00",
37544=>X"00",
37545=>X"00",
37546=>X"00",
37547=>X"00",
37548=>X"00",
37549=>X"00",
37550=>X"00",
37551=>X"00",
37552=>X"00",
37553=>X"00",
37554=>X"00",
37555=>X"00",
37556=>X"00",
37557=>X"00",
37558=>X"00",
37559=>X"00",
37560=>X"00",
37561=>X"00",
37562=>X"00",
37563=>X"00",
37564=>X"00",
37565=>X"00",
37566=>X"00",
37567=>X"00",
37568=>X"00",
37569=>X"00",
37570=>X"00",
37571=>X"00",
37572=>X"00",
37573=>X"00",
37574=>X"00",
37575=>X"00",
37576=>X"00",
37577=>X"00",
37578=>X"00",
37579=>X"00",
37580=>X"00",
37581=>X"00",
37582=>X"00",
37583=>X"00",
37584=>X"00",
37585=>X"00",
37586=>X"00",
37587=>X"00",
37588=>X"00",
37589=>X"00",
37590=>X"00",
37591=>X"00",
37592=>X"00",
37593=>X"00",
37594=>X"00",
37595=>X"00",
37596=>X"00",
37597=>X"00",
37598=>X"00",
37599=>X"00",
37600=>X"00",
37601=>X"00",
37602=>X"00",
37603=>X"00",
37604=>X"00",
37605=>X"00",
37606=>X"00",
37607=>X"00",
37608=>X"00",
37609=>X"00",
37610=>X"00",
37611=>X"00",
37612=>X"00",
37613=>X"00",
37614=>X"00",
37615=>X"00",
37616=>X"00",
37617=>X"00",
37618=>X"00",
37619=>X"00",
37620=>X"00",
37621=>X"00",
37622=>X"00",
37623=>X"00",
37624=>X"00",
37625=>X"00",
37626=>X"00",
37627=>X"00",
37628=>X"00",
37629=>X"00",
37630=>X"00",
37631=>X"00",
37632=>X"00",
37633=>X"00",
37634=>X"00",
37635=>X"00",
37636=>X"00",
37637=>X"00",
37638=>X"00",
37639=>X"00",
37640=>X"00",
37641=>X"00",
37642=>X"00",
37643=>X"00",
37644=>X"00",
37645=>X"00",
37646=>X"00",
37647=>X"00",
37648=>X"00",
37649=>X"00",
37650=>X"00",
37651=>X"00",
37652=>X"00",
37653=>X"00",
37654=>X"00",
37655=>X"00",
37656=>X"00",
37657=>X"00",
37658=>X"00",
37659=>X"00",
37660=>X"00",
37661=>X"00",
37662=>X"00",
37663=>X"00",
37664=>X"00",
37665=>X"00",
37666=>X"00",
37667=>X"00",
37668=>X"00",
37669=>X"00",
37670=>X"00",
37671=>X"00",
37672=>X"00",
37673=>X"00",
37674=>X"00",
37675=>X"00",
37676=>X"00",
37677=>X"00",
37678=>X"00",
37679=>X"00",
37680=>X"00",
37681=>X"00",
37682=>X"00",
37683=>X"00",
37684=>X"00",
37685=>X"00",
37686=>X"00",
37687=>X"00",
37688=>X"00",
37689=>X"00",
37690=>X"00",
37691=>X"00",
37692=>X"00",
37693=>X"00",
37694=>X"00",
37695=>X"00",
37696=>X"00",
37697=>X"00",
37698=>X"00",
37699=>X"00",
37700=>X"00",
37701=>X"00",
37702=>X"00",
37703=>X"00",
37704=>X"00",
37705=>X"00",
37706=>X"00",
37707=>X"00",
37708=>X"00",
37709=>X"00",
37710=>X"00",
37711=>X"00",
37712=>X"00",
37713=>X"00",
37714=>X"00",
37715=>X"00",
37716=>X"00",
37717=>X"00",
37718=>X"00",
37719=>X"00",
37720=>X"00",
37721=>X"00",
37722=>X"00",
37723=>X"00",
37724=>X"00",
37725=>X"00",
37726=>X"00",
37727=>X"00",
37728=>X"00",
37729=>X"00",
37730=>X"00",
37731=>X"00",
37732=>X"00",
37733=>X"00",
37734=>X"00",
37735=>X"00",
37736=>X"00",
37737=>X"00",
37738=>X"00",
37739=>X"00",
37740=>X"00",
37741=>X"00",
37742=>X"00",
37743=>X"00",
37744=>X"00",
37745=>X"00",
37746=>X"00",
37747=>X"00",
37748=>X"00",
37749=>X"00",
37750=>X"00",
37751=>X"00",
37752=>X"00",
37753=>X"00",
37754=>X"00",
37755=>X"00",
37756=>X"00",
37757=>X"00",
37758=>X"00",
37759=>X"00",
37760=>X"00",
37761=>X"00",
37762=>X"00",
37763=>X"00",
37764=>X"00",
37765=>X"00",
37766=>X"00",
37767=>X"00",
37768=>X"00",
37769=>X"00",
37770=>X"00",
37771=>X"00",
37772=>X"00",
37773=>X"00",
37774=>X"00",
37775=>X"00",
37776=>X"00",
37777=>X"00",
37778=>X"00",
37779=>X"00",
37780=>X"00",
37781=>X"00",
37782=>X"00",
37783=>X"00",
37784=>X"00",
37785=>X"00",
37786=>X"00",
37787=>X"00",
37788=>X"00",
37789=>X"00",
37790=>X"00",
37791=>X"00",
37792=>X"00",
37793=>X"00",
37794=>X"00",
37795=>X"00",
37796=>X"00",
37797=>X"00",
37798=>X"00",
37799=>X"00",
37800=>X"00",
37801=>X"00",
37802=>X"00",
37803=>X"00",
37804=>X"00",
37805=>X"00",
37806=>X"00",
37807=>X"00",
37808=>X"00",
37809=>X"00",
37810=>X"00",
37811=>X"00",
37812=>X"00",
37813=>X"00",
37814=>X"00",
37815=>X"00",
37816=>X"00",
37817=>X"00",
37818=>X"00",
37819=>X"00",
37820=>X"00",
37821=>X"00",
37822=>X"00",
37823=>X"00",
37824=>X"00",
37825=>X"00",
37826=>X"00",
37827=>X"00",
37828=>X"00",
37829=>X"00",
37830=>X"00",
37831=>X"00",
37832=>X"00",
37833=>X"00",
37834=>X"00",
37835=>X"00",
37836=>X"00",
37837=>X"00",
37838=>X"00",
37839=>X"00",
37840=>X"00",
37841=>X"00",
37842=>X"00",
37843=>X"00",
37844=>X"00",
37845=>X"00",
37846=>X"00",
37847=>X"00",
37848=>X"00",
37849=>X"00",
37850=>X"00",
37851=>X"00",
37852=>X"00",
37853=>X"00",
37854=>X"00",
37855=>X"00",
37856=>X"00",
37857=>X"00",
37858=>X"00",
37859=>X"00",
37860=>X"00",
37861=>X"00",
37862=>X"00",
37863=>X"00",
37864=>X"00",
37865=>X"00",
37866=>X"00",
37867=>X"00",
37868=>X"00",
37869=>X"00",
37870=>X"00",
37871=>X"00",
37872=>X"00",
37873=>X"00",
37874=>X"00",
37875=>X"00",
37876=>X"00",
37877=>X"00",
37878=>X"00",
37879=>X"00",
37880=>X"00",
37881=>X"00",
37882=>X"00",
37883=>X"00",
37884=>X"00",
37885=>X"00",
37886=>X"00",
37887=>X"00",
37888=>X"00",
37889=>X"00",
37890=>X"00",
37891=>X"00",
37892=>X"00",
37893=>X"00",
37894=>X"00",
37895=>X"00",
37896=>X"00",
37897=>X"00",
37898=>X"00",
37899=>X"00",
37900=>X"00",
37901=>X"00",
37902=>X"00",
37903=>X"00",
37904=>X"00",
37905=>X"00",
37906=>X"00",
37907=>X"00",
37908=>X"00",
37909=>X"00",
37910=>X"00",
37911=>X"00",
37912=>X"00",
37913=>X"00",
37914=>X"00",
37915=>X"00",
37916=>X"00",
37917=>X"00",
37918=>X"00",
37919=>X"00",
37920=>X"00",
37921=>X"00",
37922=>X"00",
37923=>X"00",
37924=>X"00",
37925=>X"00",
37926=>X"00",
37927=>X"00",
37928=>X"00",
37929=>X"00",
37930=>X"00",
37931=>X"00",
37932=>X"00",
37933=>X"00",
37934=>X"00",
37935=>X"00",
37936=>X"00",
37937=>X"00",
37938=>X"00",
37939=>X"00",
37940=>X"00",
37941=>X"00",
37942=>X"00",
37943=>X"00",
37944=>X"00",
37945=>X"00",
37946=>X"00",
37947=>X"00",
37948=>X"00",
37949=>X"00",
37950=>X"00",
37951=>X"00",
37952=>X"00",
37953=>X"00",
37954=>X"00",
37955=>X"00",
37956=>X"00",
37957=>X"00",
37958=>X"00",
37959=>X"00",
37960=>X"00",
37961=>X"00",
37962=>X"00",
37963=>X"00",
37964=>X"00",
37965=>X"00",
37966=>X"00",
37967=>X"00",
37968=>X"00",
37969=>X"00",
37970=>X"00",
37971=>X"00",
37972=>X"00",
37973=>X"00",
37974=>X"00",
37975=>X"00",
37976=>X"00",
37977=>X"00",
37978=>X"00",
37979=>X"00",
37980=>X"00",
37981=>X"00",
37982=>X"00",
37983=>X"00",
37984=>X"00",
37985=>X"00",
37986=>X"00",
37987=>X"00",
37988=>X"00",
37989=>X"00",
37990=>X"00",
37991=>X"00",
37992=>X"00",
37993=>X"00",
37994=>X"00",
37995=>X"00",
37996=>X"00",
37997=>X"00",
37998=>X"00",
37999=>X"00",
38000=>X"00",
38001=>X"00",
38002=>X"00",
38003=>X"00",
38004=>X"00",
38005=>X"00",
38006=>X"00",
38007=>X"00",
38008=>X"00",
38009=>X"00",
38010=>X"00",
38011=>X"00",
38012=>X"00",
38013=>X"00",
38014=>X"00",
38015=>X"00",
38016=>X"00",
38017=>X"00",
38018=>X"00",
38019=>X"00",
38020=>X"00",
38021=>X"00",
38022=>X"00",
38023=>X"00",
38024=>X"00",
38025=>X"00",
38026=>X"00",
38027=>X"00",
38028=>X"00",
38029=>X"00",
38030=>X"00",
38031=>X"00",
38032=>X"00",
38033=>X"00",
38034=>X"00",
38035=>X"00",
38036=>X"00",
38037=>X"00",
38038=>X"00",
38039=>X"00",
38040=>X"00",
38041=>X"00",
38042=>X"00",
38043=>X"00",
38044=>X"00",
38045=>X"00",
38046=>X"00",
38047=>X"00",
38048=>X"00",
38049=>X"00",
38050=>X"00",
38051=>X"00",
38052=>X"00",
38053=>X"00",
38054=>X"00",
38055=>X"00",
38056=>X"00",
38057=>X"00",
38058=>X"00",
38059=>X"00",
38060=>X"00",
38061=>X"00",
38062=>X"00",
38063=>X"00",
38064=>X"00",
38065=>X"00",
38066=>X"00",
38067=>X"00",
38068=>X"00",
38069=>X"00",
38070=>X"00",
38071=>X"00",
38072=>X"00",
38073=>X"00",
38074=>X"00",
38075=>X"00",
38076=>X"00",
38077=>X"00",
38078=>X"00",
38079=>X"00",
38080=>X"00",
38081=>X"00",
38082=>X"00",
38083=>X"00",
38084=>X"00",
38085=>X"00",
38086=>X"00",
38087=>X"00",
38088=>X"00",
38089=>X"00",
38090=>X"00",
38091=>X"00",
38092=>X"00",
38093=>X"00",
38094=>X"00",
38095=>X"00",
38096=>X"00",
38097=>X"00",
38098=>X"00",
38099=>X"00",
38100=>X"00",
38101=>X"00",
38102=>X"00",
38103=>X"00",
38104=>X"00",
38105=>X"00",
38106=>X"00",
38107=>X"00",
38108=>X"00",
38109=>X"00",
38110=>X"00",
38111=>X"00",
38112=>X"00",
38113=>X"00",
38114=>X"00",
38115=>X"00",
38116=>X"00",
38117=>X"00",
38118=>X"00",
38119=>X"00",
38120=>X"00",
38121=>X"00",
38122=>X"00",
38123=>X"00",
38124=>X"00",
38125=>X"00",
38126=>X"00",
38127=>X"00",
38128=>X"00",
38129=>X"00",
38130=>X"00",
38131=>X"00",
38132=>X"00",
38133=>X"00",
38134=>X"00",
38135=>X"00",
38136=>X"00",
38137=>X"00",
38138=>X"00",
38139=>X"00",
38140=>X"00",
38141=>X"00",
38142=>X"00",
38143=>X"00",
38144=>X"00",
38145=>X"00",
38146=>X"00",
38147=>X"00",
38148=>X"00",
38149=>X"00",
38150=>X"00",
38151=>X"00",
38152=>X"00",
38153=>X"00",
38154=>X"00",
38155=>X"00",
38156=>X"00",
38157=>X"00",
38158=>X"00",
38159=>X"00",
38160=>X"00",
38161=>X"00",
38162=>X"00",
38163=>X"00",
38164=>X"00",
38165=>X"00",
38166=>X"00",
38167=>X"00",
38168=>X"00",
38169=>X"00",
38170=>X"00",
38171=>X"00",
38172=>X"00",
38173=>X"00",
38174=>X"00",
38175=>X"00",
38176=>X"00",
38177=>X"00",
38178=>X"00",
38179=>X"00",
38180=>X"00",
38181=>X"00",
38182=>X"00",
38183=>X"00",
38184=>X"00",
38185=>X"00",
38186=>X"00",
38187=>X"00",
38188=>X"00",
38189=>X"00",
38190=>X"00",
38191=>X"00",
38192=>X"00",
38193=>X"00",
38194=>X"00",
38195=>X"00",
38196=>X"00",
38197=>X"00",
38198=>X"00",
38199=>X"00",
38200=>X"00",
38201=>X"00",
38202=>X"00",
38203=>X"00",
38204=>X"00",
38205=>X"00",
38206=>X"00",
38207=>X"00",
38208=>X"00",
38209=>X"00",
38210=>X"00",
38211=>X"00",
38212=>X"00",
38213=>X"00",
38214=>X"00",
38215=>X"00",
38216=>X"00",
38217=>X"00",
38218=>X"00",
38219=>X"00",
38220=>X"00",
38221=>X"00",
38222=>X"00",
38223=>X"00",
38224=>X"00",
38225=>X"00",
38226=>X"00",
38227=>X"00",
38228=>X"00",
38229=>X"00",
38230=>X"00",
38231=>X"00",
38232=>X"00",
38233=>X"00",
38234=>X"00",
38235=>X"00",
38236=>X"00",
38237=>X"00",
38238=>X"00",
38239=>X"00",
38240=>X"00",
38241=>X"00",
38242=>X"00",
38243=>X"00",
38244=>X"00",
38245=>X"00",
38246=>X"00",
38247=>X"00",
38248=>X"00",
38249=>X"00",
38250=>X"00",
38251=>X"00",
38252=>X"00",
38253=>X"00",
38254=>X"00",
38255=>X"00",
38256=>X"00",
38257=>X"00",
38258=>X"00",
38259=>X"00",
38260=>X"00",
38261=>X"00",
38262=>X"00",
38263=>X"00",
38264=>X"00",
38265=>X"00",
38266=>X"00",
38267=>X"00",
38268=>X"00",
38269=>X"00",
38270=>X"00",
38271=>X"00",
38272=>X"00",
38273=>X"00",
38274=>X"00",
38275=>X"00",
38276=>X"00",
38277=>X"00",
38278=>X"00",
38279=>X"00",
38280=>X"00",
38281=>X"00",
38282=>X"00",
38283=>X"00",
38284=>X"00",
38285=>X"00",
38286=>X"00",
38287=>X"00",
38288=>X"00",
38289=>X"00",
38290=>X"00",
38291=>X"00",
38292=>X"00",
38293=>X"00",
38294=>X"00",
38295=>X"00",
38296=>X"00",
38297=>X"00",
38298=>X"00",
38299=>X"00",
38300=>X"00",
38301=>X"00",
38302=>X"00",
38303=>X"00",
38304=>X"00",
38305=>X"00",
38306=>X"00",
38307=>X"00",
38308=>X"00",
38309=>X"00",
38310=>X"00",
38311=>X"00",
38312=>X"00",
38313=>X"00",
38314=>X"00",
38315=>X"00",
38316=>X"00",
38317=>X"00",
38318=>X"00",
38319=>X"00",
38320=>X"00",
38321=>X"00",
38322=>X"00",
38323=>X"00",
38324=>X"00",
38325=>X"00",
38326=>X"00",
38327=>X"00",
38328=>X"00",
38329=>X"00",
38330=>X"00",
38331=>X"00",
38332=>X"00",
38333=>X"00",
38334=>X"00",
38335=>X"00",
38336=>X"00",
38337=>X"00",
38338=>X"00",
38339=>X"00",
38340=>X"00",
38341=>X"00",
38342=>X"00",
38343=>X"00",
38344=>X"00",
38345=>X"00",
38346=>X"00",
38347=>X"00",
38348=>X"00",
38349=>X"00",
38350=>X"00",
38351=>X"00",
38352=>X"00",
38353=>X"00",
38354=>X"00",
38355=>X"00",
38356=>X"00",
38357=>X"00",
38358=>X"00",
38359=>X"00",
38360=>X"00",
38361=>X"00",
38362=>X"00",
38363=>X"00",
38364=>X"00",
38365=>X"00",
38366=>X"00",
38367=>X"00",
38368=>X"00",
38369=>X"00",
38370=>X"00",
38371=>X"00",
38372=>X"00",
38373=>X"00",
38374=>X"00",
38375=>X"00",
38376=>X"00",
38377=>X"00",
38378=>X"00",
38379=>X"00",
38380=>X"00",
38381=>X"00",
38382=>X"00",
38383=>X"00",
38384=>X"00",
38385=>X"00",
38386=>X"00",
38387=>X"00",
38388=>X"00",
38389=>X"00",
38390=>X"00",
38391=>X"00",
38392=>X"00",
38393=>X"00",
38394=>X"00",
38395=>X"00",
38396=>X"00",
38397=>X"00",
38398=>X"00",
38399=>X"00",
38400=>X"00",
38401=>X"00",
38402=>X"00",
38403=>X"00",
38404=>X"00",
38405=>X"00",
38406=>X"00",
38407=>X"00",
38408=>X"00",
38409=>X"00",
38410=>X"00",
38411=>X"00",
38412=>X"00",
38413=>X"00",
38414=>X"00",
38415=>X"00",
38416=>X"00",
38417=>X"00",
38418=>X"00",
38419=>X"00",
38420=>X"00",
38421=>X"00",
38422=>X"00",
38423=>X"00",
38424=>X"00",
38425=>X"00",
38426=>X"00",
38427=>X"00",
38428=>X"00",
38429=>X"00",
38430=>X"00",
38431=>X"00",
38432=>X"00",
38433=>X"00",
38434=>X"00",
38435=>X"00",
38436=>X"00",
38437=>X"00",
38438=>X"00",
38439=>X"00",
38440=>X"00",
38441=>X"00",
38442=>X"00",
38443=>X"00",
38444=>X"00",
38445=>X"00",
38446=>X"00",
38447=>X"00",
38448=>X"00",
38449=>X"00",
38450=>X"00",
38451=>X"00",
38452=>X"00",
38453=>X"00",
38454=>X"00",
38455=>X"00",
38456=>X"00",
38457=>X"00",
38458=>X"00",
38459=>X"00",
38460=>X"00",
38461=>X"00",
38462=>X"00",
38463=>X"00",
38464=>X"00",
38465=>X"00",
38466=>X"00",
38467=>X"00",
38468=>X"00",
38469=>X"00",
38470=>X"00",
38471=>X"00",
38472=>X"00",
38473=>X"00",
38474=>X"00",
38475=>X"00",
38476=>X"00",
38477=>X"00",
38478=>X"00",
38479=>X"00",
38480=>X"00",
38481=>X"00",
38482=>X"00",
38483=>X"00",
38484=>X"00",
38485=>X"00",
38486=>X"00",
38487=>X"00",
38488=>X"00",
38489=>X"00",
38490=>X"00",
38491=>X"00",
38492=>X"00",
38493=>X"00",
38494=>X"00",
38495=>X"00",
38496=>X"00",
38497=>X"00",
38498=>X"00",
38499=>X"00",
38500=>X"00",
38501=>X"00",
38502=>X"00",
38503=>X"00",
38504=>X"00",
38505=>X"00",
38506=>X"00",
38507=>X"00",
38508=>X"00",
38509=>X"00",
38510=>X"00",
38511=>X"00",
38512=>X"00",
38513=>X"00",
38514=>X"00",
38515=>X"00",
38516=>X"00",
38517=>X"00",
38518=>X"00",
38519=>X"00",
38520=>X"00",
38521=>X"00",
38522=>X"00",
38523=>X"00",
38524=>X"00",
38525=>X"00",
38526=>X"00",
38527=>X"00",
38528=>X"00",
38529=>X"00",
38530=>X"00",
38531=>X"00",
38532=>X"00",
38533=>X"00",
38534=>X"00",
38535=>X"00",
38536=>X"00",
38537=>X"00",
38538=>X"00",
38539=>X"00",
38540=>X"00",
38541=>X"00",
38542=>X"00",
38543=>X"00",
38544=>X"00",
38545=>X"00",
38546=>X"00",
38547=>X"00",
38548=>X"00",
38549=>X"00",
38550=>X"00",
38551=>X"00",
38552=>X"00",
38553=>X"00",
38554=>X"00",
38555=>X"00",
38556=>X"00",
38557=>X"00",
38558=>X"00",
38559=>X"00",
38560=>X"00",
38561=>X"00",
38562=>X"00",
38563=>X"00",
38564=>X"00",
38565=>X"00",
38566=>X"00",
38567=>X"00",
38568=>X"00",
38569=>X"00",
38570=>X"00",
38571=>X"00",
38572=>X"00",
38573=>X"00",
38574=>X"00",
38575=>X"00",
38576=>X"00",
38577=>X"00",
38578=>X"00",
38579=>X"00",
38580=>X"00",
38581=>X"00",
38582=>X"00",
38583=>X"00",
38584=>X"00",
38585=>X"00",
38586=>X"00",
38587=>X"00",
38588=>X"00",
38589=>X"00",
38590=>X"00",
38591=>X"00",
38592=>X"00",
38593=>X"00",
38594=>X"00",
38595=>X"00",
38596=>X"00",
38597=>X"00",
38598=>X"00",
38599=>X"00",
38600=>X"00",
38601=>X"00",
38602=>X"00",
38603=>X"00",
38604=>X"00",
38605=>X"00",
38606=>X"00",
38607=>X"00",
38608=>X"00",
38609=>X"00",
38610=>X"00",
38611=>X"00",
38612=>X"00",
38613=>X"00",
38614=>X"00",
38615=>X"00",
38616=>X"00",
38617=>X"00",
38618=>X"00",
38619=>X"00",
38620=>X"00",
38621=>X"00",
38622=>X"00",
38623=>X"00",
38624=>X"00",
38625=>X"00",
38626=>X"00",
38627=>X"00",
38628=>X"00",
38629=>X"00",
38630=>X"00",
38631=>X"00",
38632=>X"00",
38633=>X"00",
38634=>X"00",
38635=>X"00",
38636=>X"00",
38637=>X"00",
38638=>X"00",
38639=>X"00",
38640=>X"00",
38641=>X"00",
38642=>X"00",
38643=>X"00",
38644=>X"00",
38645=>X"00",
38646=>X"00",
38647=>X"00",
38648=>X"00",
38649=>X"00",
38650=>X"00",
38651=>X"00",
38652=>X"00",
38653=>X"00",
38654=>X"00",
38655=>X"00",
38656=>X"00",
38657=>X"00",
38658=>X"00",
38659=>X"00",
38660=>X"00",
38661=>X"00",
38662=>X"00",
38663=>X"00",
38664=>X"00",
38665=>X"00",
38666=>X"00",
38667=>X"00",
38668=>X"00",
38669=>X"00",
38670=>X"00",
38671=>X"00",
38672=>X"00",
38673=>X"00",
38674=>X"00",
38675=>X"00",
38676=>X"00",
38677=>X"00",
38678=>X"00",
38679=>X"00",
38680=>X"00",
38681=>X"00",
38682=>X"00",
38683=>X"00",
38684=>X"00",
38685=>X"00",
38686=>X"00",
38687=>X"00",
38688=>X"00",
38689=>X"00",
38690=>X"00",
38691=>X"00",
38692=>X"00",
38693=>X"00",
38694=>X"00",
38695=>X"00",
38696=>X"00",
38697=>X"00",
38698=>X"00",
38699=>X"00",
38700=>X"00",
38701=>X"00",
38702=>X"00",
38703=>X"00",
38704=>X"00",
38705=>X"00",
38706=>X"00",
38707=>X"00",
38708=>X"00",
38709=>X"00",
38710=>X"00",
38711=>X"00",
38712=>X"00",
38713=>X"00",
38714=>X"00",
38715=>X"00",
38716=>X"00",
38717=>X"00",
38718=>X"00",
38719=>X"00",
38720=>X"00",
38721=>X"00",
38722=>X"00",
38723=>X"00",
38724=>X"00",
38725=>X"00",
38726=>X"00",
38727=>X"00",
38728=>X"00",
38729=>X"00",
38730=>X"00",
38731=>X"00",
38732=>X"00",
38733=>X"00",
38734=>X"00",
38735=>X"00",
38736=>X"00",
38737=>X"00",
38738=>X"00",
38739=>X"00",
38740=>X"00",
38741=>X"00",
38742=>X"00",
38743=>X"00",
38744=>X"00",
38745=>X"00",
38746=>X"00",
38747=>X"00",
38748=>X"00",
38749=>X"00",
38750=>X"00",
38751=>X"00",
38752=>X"00",
38753=>X"00",
38754=>X"00",
38755=>X"00",
38756=>X"00",
38757=>X"00",
38758=>X"00",
38759=>X"00",
38760=>X"00",
38761=>X"00",
38762=>X"00",
38763=>X"00",
38764=>X"00",
38765=>X"00",
38766=>X"00",
38767=>X"00",
38768=>X"00",
38769=>X"00",
38770=>X"00",
38771=>X"00",
38772=>X"00",
38773=>X"00",
38774=>X"00",
38775=>X"00",
38776=>X"00",
38777=>X"00",
38778=>X"00",
38779=>X"00",
38780=>X"00",
38781=>X"00",
38782=>X"00",
38783=>X"00",
38784=>X"00",
38785=>X"00",
38786=>X"00",
38787=>X"00",
38788=>X"00",
38789=>X"00",
38790=>X"00",
38791=>X"00",
38792=>X"00",
38793=>X"00",
38794=>X"00",
38795=>X"00",
38796=>X"00",
38797=>X"00",
38798=>X"00",
38799=>X"00",
38800=>X"00",
38801=>X"00",
38802=>X"00",
38803=>X"00",
38804=>X"00",
38805=>X"00",
38806=>X"00",
38807=>X"00",
38808=>X"00",
38809=>X"00",
38810=>X"00",
38811=>X"00",
38812=>X"00",
38813=>X"00",
38814=>X"00",
38815=>X"00",
38816=>X"00",
38817=>X"00",
38818=>X"00",
38819=>X"00",
38820=>X"00",
38821=>X"00",
38822=>X"00",
38823=>X"00",
38824=>X"00",
38825=>X"00",
38826=>X"00",
38827=>X"00",
38828=>X"00",
38829=>X"00",
38830=>X"00",
38831=>X"00",
38832=>X"00",
38833=>X"00",
38834=>X"00",
38835=>X"00",
38836=>X"00",
38837=>X"00",
38838=>X"00",
38839=>X"00",
38840=>X"00",
38841=>X"00",
38842=>X"00",
38843=>X"00",
38844=>X"00",
38845=>X"00",
38846=>X"00",
38847=>X"00",
38848=>X"00",
38849=>X"00",
38850=>X"00",
38851=>X"00",
38852=>X"00",
38853=>X"00",
38854=>X"00",
38855=>X"00",
38856=>X"00",
38857=>X"00",
38858=>X"00",
38859=>X"00",
38860=>X"00",
38861=>X"00",
38862=>X"00",
38863=>X"00",
38864=>X"00",
38865=>X"00",
38866=>X"00",
38867=>X"00",
38868=>X"00",
38869=>X"00",
38870=>X"00",
38871=>X"00",
38872=>X"00",
38873=>X"00",
38874=>X"00",
38875=>X"00",
38876=>X"00",
38877=>X"00",
38878=>X"00",
38879=>X"00",
38880=>X"00",
38881=>X"00",
38882=>X"00",
38883=>X"00",
38884=>X"00",
38885=>X"00",
38886=>X"00",
38887=>X"00",
38888=>X"00",
38889=>X"00",
38890=>X"00",
38891=>X"00",
38892=>X"00",
38893=>X"00",
38894=>X"00",
38895=>X"00",
38896=>X"00",
38897=>X"00",
38898=>X"00",
38899=>X"00",
38900=>X"00",
38901=>X"00",
38902=>X"00",
38903=>X"00",
38904=>X"00",
38905=>X"00",
38906=>X"00",
38907=>X"00",
38908=>X"00",
38909=>X"00",
38910=>X"00",
38911=>X"00",
38912=>X"00",
38913=>X"00",
38914=>X"00",
38915=>X"00",
38916=>X"00",
38917=>X"00",
38918=>X"00",
38919=>X"00",
38920=>X"00",
38921=>X"00",
38922=>X"00",
38923=>X"00",
38924=>X"00",
38925=>X"00",
38926=>X"00",
38927=>X"00",
38928=>X"00",
38929=>X"00",
38930=>X"00",
38931=>X"00",
38932=>X"00",
38933=>X"00",
38934=>X"00",
38935=>X"00",
38936=>X"00",
38937=>X"00",
38938=>X"00",
38939=>X"00",
38940=>X"00",
38941=>X"00",
38942=>X"00",
38943=>X"00",
38944=>X"00",
38945=>X"00",
38946=>X"00",
38947=>X"00",
38948=>X"00",
38949=>X"00",
38950=>X"00",
38951=>X"00",
38952=>X"00",
38953=>X"00",
38954=>X"00",
38955=>X"00",
38956=>X"00",
38957=>X"00",
38958=>X"00",
38959=>X"00",
38960=>X"00",
38961=>X"00",
38962=>X"00",
38963=>X"00",
38964=>X"00",
38965=>X"00",
38966=>X"00",
38967=>X"00",
38968=>X"00",
38969=>X"00",
38970=>X"00",
38971=>X"00",
38972=>X"00",
38973=>X"00",
38974=>X"00",
38975=>X"00",
38976=>X"00",
38977=>X"00",
38978=>X"00",
38979=>X"00",
38980=>X"00",
38981=>X"00",
38982=>X"00",
38983=>X"00",
38984=>X"00",
38985=>X"00",
38986=>X"00",
38987=>X"00",
38988=>X"00",
38989=>X"00",
38990=>X"00",
38991=>X"00",
38992=>X"00",
38993=>X"00",
38994=>X"00",
38995=>X"00",
38996=>X"00",
38997=>X"00",
38998=>X"00",
38999=>X"00",
39000=>X"00",
39001=>X"00",
39002=>X"00",
39003=>X"00",
39004=>X"00",
39005=>X"00",
39006=>X"00",
39007=>X"00",
39008=>X"00",
39009=>X"00",
39010=>X"00",
39011=>X"00",
39012=>X"00",
39013=>X"00",
39014=>X"00",
39015=>X"00",
39016=>X"00",
39017=>X"00",
39018=>X"00",
39019=>X"00",
39020=>X"00",
39021=>X"00",
39022=>X"00",
39023=>X"00",
39024=>X"00",
39025=>X"00",
39026=>X"00",
39027=>X"00",
39028=>X"00",
39029=>X"00",
39030=>X"00",
39031=>X"00",
39032=>X"00",
39033=>X"00",
39034=>X"00",
39035=>X"00",
39036=>X"00",
39037=>X"00",
39038=>X"00",
39039=>X"00",
39040=>X"00",
39041=>X"00",
39042=>X"00",
39043=>X"00",
39044=>X"00",
39045=>X"00",
39046=>X"00",
39047=>X"00",
39048=>X"00",
39049=>X"00",
39050=>X"00",
39051=>X"00",
39052=>X"00",
39053=>X"00",
39054=>X"00",
39055=>X"00",
39056=>X"00",
39057=>X"00",
39058=>X"00",
39059=>X"00",
39060=>X"00",
39061=>X"00",
39062=>X"00",
39063=>X"00",
39064=>X"00",
39065=>X"00",
39066=>X"00",
39067=>X"00",
39068=>X"00",
39069=>X"00",
39070=>X"00",
39071=>X"00",
39072=>X"00",
39073=>X"00",
39074=>X"00",
39075=>X"00",
39076=>X"00",
39077=>X"00",
39078=>X"00",
39079=>X"00",
39080=>X"00",
39081=>X"00",
39082=>X"00",
39083=>X"00",
39084=>X"00",
39085=>X"00",
39086=>X"00",
39087=>X"00",
39088=>X"00",
39089=>X"00",
39090=>X"00",
39091=>X"00",
39092=>X"00",
39093=>X"00",
39094=>X"00",
39095=>X"00",
39096=>X"00",
39097=>X"00",
39098=>X"00",
39099=>X"00",
39100=>X"00",
39101=>X"00",
39102=>X"00",
39103=>X"00",
39104=>X"00",
39105=>X"00",
39106=>X"00",
39107=>X"00",
39108=>X"00",
39109=>X"00",
39110=>X"00",
39111=>X"00",
39112=>X"00",
39113=>X"00",
39114=>X"00",
39115=>X"00",
39116=>X"00",
39117=>X"00",
39118=>X"00",
39119=>X"00",
39120=>X"00",
39121=>X"00",
39122=>X"00",
39123=>X"00",
39124=>X"00",
39125=>X"00",
39126=>X"00",
39127=>X"00",
39128=>X"00",
39129=>X"00",
39130=>X"00",
39131=>X"00",
39132=>X"00",
39133=>X"00",
39134=>X"00",
39135=>X"00",
39136=>X"00",
39137=>X"00",
39138=>X"00",
39139=>X"00",
39140=>X"00",
39141=>X"00",
39142=>X"00",
39143=>X"00",
39144=>X"00",
39145=>X"00",
39146=>X"00",
39147=>X"00",
39148=>X"00",
39149=>X"00",
39150=>X"00",
39151=>X"00",
39152=>X"00",
39153=>X"00",
39154=>X"00",
39155=>X"00",
39156=>X"00",
39157=>X"00",
39158=>X"00",
39159=>X"00",
39160=>X"00",
39161=>X"00",
39162=>X"00",
39163=>X"00",
39164=>X"00",
39165=>X"00",
39166=>X"00",
39167=>X"00",
39168=>X"00",
39169=>X"00",
39170=>X"00",
39171=>X"00",
39172=>X"00",
39173=>X"00",
39174=>X"00",
39175=>X"00",
39176=>X"00",
39177=>X"00",
39178=>X"00",
39179=>X"00",
39180=>X"00",
39181=>X"00",
39182=>X"00",
39183=>X"00",
39184=>X"00",
39185=>X"00",
39186=>X"00",
39187=>X"00",
39188=>X"00",
39189=>X"00",
39190=>X"00",
39191=>X"00",
39192=>X"00",
39193=>X"00",
39194=>X"00",
39195=>X"00",
39196=>X"00",
39197=>X"00",
39198=>X"00",
39199=>X"00",
39200=>X"00",
39201=>X"00",
39202=>X"00",
39203=>X"00",
39204=>X"00",
39205=>X"00",
39206=>X"00",
39207=>X"00",
39208=>X"00",
39209=>X"00",
39210=>X"00",
39211=>X"00",
39212=>X"00",
39213=>X"00",
39214=>X"00",
39215=>X"00",
39216=>X"00",
39217=>X"00",
39218=>X"00",
39219=>X"00",
39220=>X"00",
39221=>X"00",
39222=>X"00",
39223=>X"00",
39224=>X"00",
39225=>X"00",
39226=>X"00",
39227=>X"00",
39228=>X"00",
39229=>X"00",
39230=>X"00",
39231=>X"00",
39232=>X"00",
39233=>X"00",
39234=>X"00",
39235=>X"00",
39236=>X"00",
39237=>X"00",
39238=>X"00",
39239=>X"00",
39240=>X"00",
39241=>X"00",
39242=>X"00",
39243=>X"00",
39244=>X"00",
39245=>X"00",
39246=>X"00",
39247=>X"00",
39248=>X"00",
39249=>X"00",
39250=>X"00",
39251=>X"00",
39252=>X"00",
39253=>X"00",
39254=>X"00",
39255=>X"00",
39256=>X"00",
39257=>X"00",
39258=>X"00",
39259=>X"00",
39260=>X"00",
39261=>X"00",
39262=>X"00",
39263=>X"00",
39264=>X"00",
39265=>X"00",
39266=>X"00",
39267=>X"00",
39268=>X"00",
39269=>X"00",
39270=>X"00",
39271=>X"00",
39272=>X"00",
39273=>X"00",
39274=>X"00",
39275=>X"00",
39276=>X"00",
39277=>X"00",
39278=>X"00",
39279=>X"00",
39280=>X"00",
39281=>X"00",
39282=>X"00",
39283=>X"00",
39284=>X"00",
39285=>X"00",
39286=>X"00",
39287=>X"00",
39288=>X"00",
39289=>X"00",
39290=>X"00",
39291=>X"00",
39292=>X"00",
39293=>X"00",
39294=>X"00",
39295=>X"00",
39296=>X"00",
39297=>X"00",
39298=>X"00",
39299=>X"00",
39300=>X"00",
39301=>X"00",
39302=>X"00",
39303=>X"00",
39304=>X"00",
39305=>X"00",
39306=>X"00",
39307=>X"00",
39308=>X"00",
39309=>X"00",
39310=>X"00",
39311=>X"00",
39312=>X"00",
39313=>X"00",
39314=>X"00",
39315=>X"00",
39316=>X"00",
39317=>X"00",
39318=>X"00",
39319=>X"00",
39320=>X"00",
39321=>X"00",
39322=>X"00",
39323=>X"00",
39324=>X"00",
39325=>X"00",
39326=>X"00",
39327=>X"00",
39328=>X"00",
39329=>X"00",
39330=>X"00",
39331=>X"00",
39332=>X"00",
39333=>X"00",
39334=>X"00",
39335=>X"00",
39336=>X"00",
39337=>X"00",
39338=>X"00",
39339=>X"00",
39340=>X"00",
39341=>X"00",
39342=>X"00",
39343=>X"00",
39344=>X"00",
39345=>X"00",
39346=>X"00",
39347=>X"00",
39348=>X"00",
39349=>X"00",
39350=>X"00",
39351=>X"00",
39352=>X"00",
39353=>X"00",
39354=>X"00",
39355=>X"00",
39356=>X"00",
39357=>X"00",
39358=>X"00",
39359=>X"00",
39360=>X"00",
39361=>X"00",
39362=>X"00",
39363=>X"00",
39364=>X"00",
39365=>X"00",
39366=>X"00",
39367=>X"00",
39368=>X"00",
39369=>X"00",
39370=>X"00",
39371=>X"00",
39372=>X"00",
39373=>X"00",
39374=>X"00",
39375=>X"00",
39376=>X"00",
39377=>X"00",
39378=>X"00",
39379=>X"00",
39380=>X"00",
39381=>X"00",
39382=>X"00",
39383=>X"00",
39384=>X"00",
39385=>X"00",
39386=>X"00",
39387=>X"00",
39388=>X"00",
39389=>X"00",
39390=>X"00",
39391=>X"00",
39392=>X"00",
39393=>X"00",
39394=>X"00",
39395=>X"00",
39396=>X"00",
39397=>X"00",
39398=>X"00",
39399=>X"00",
39400=>X"00",
39401=>X"00",
39402=>X"00",
39403=>X"00",
39404=>X"00",
39405=>X"00",
39406=>X"00",
39407=>X"00",
39408=>X"00",
39409=>X"00",
39410=>X"00",
39411=>X"00",
39412=>X"00",
39413=>X"00",
39414=>X"00",
39415=>X"00",
39416=>X"00",
39417=>X"00",
39418=>X"00",
39419=>X"00",
39420=>X"00",
39421=>X"00",
39422=>X"00",
39423=>X"00",
39424=>X"00",
39425=>X"00",
39426=>X"00",
39427=>X"00",
39428=>X"00",
39429=>X"00",
39430=>X"00",
39431=>X"00",
39432=>X"00",
39433=>X"00",
39434=>X"00",
39435=>X"00",
39436=>X"00",
39437=>X"00",
39438=>X"00",
39439=>X"00",
39440=>X"00",
39441=>X"00",
39442=>X"00",
39443=>X"00",
39444=>X"00",
39445=>X"00",
39446=>X"00",
39447=>X"00",
39448=>X"00",
39449=>X"00",
39450=>X"00",
39451=>X"00",
39452=>X"00",
39453=>X"00",
39454=>X"00",
39455=>X"00",
39456=>X"00",
39457=>X"00",
39458=>X"00",
39459=>X"00",
39460=>X"00",
39461=>X"00",
39462=>X"00",
39463=>X"00",
39464=>X"00",
39465=>X"00",
39466=>X"00",
39467=>X"00",
39468=>X"00",
39469=>X"00",
39470=>X"00",
39471=>X"00",
39472=>X"00",
39473=>X"00",
39474=>X"00",
39475=>X"00",
39476=>X"00",
39477=>X"00",
39478=>X"00",
39479=>X"00",
39480=>X"00",
39481=>X"00",
39482=>X"00",
39483=>X"00",
39484=>X"00",
39485=>X"00",
39486=>X"00",
39487=>X"00",
39488=>X"00",
39489=>X"00",
39490=>X"00",
39491=>X"00",
39492=>X"00",
39493=>X"00",
39494=>X"00",
39495=>X"00",
39496=>X"00",
39497=>X"00",
39498=>X"00",
39499=>X"00",
39500=>X"00",
39501=>X"00",
39502=>X"00",
39503=>X"00",
39504=>X"00",
39505=>X"00",
39506=>X"00",
39507=>X"00",
39508=>X"00",
39509=>X"00",
39510=>X"00",
39511=>X"00",
39512=>X"00",
39513=>X"00",
39514=>X"00",
39515=>X"00",
39516=>X"00",
39517=>X"00",
39518=>X"00",
39519=>X"00",
39520=>X"00",
39521=>X"00",
39522=>X"00",
39523=>X"00",
39524=>X"00",
39525=>X"00",
39526=>X"00",
39527=>X"00",
39528=>X"00",
39529=>X"00",
39530=>X"00",
39531=>X"00",
39532=>X"00",
39533=>X"00",
39534=>X"00",
39535=>X"00",
39536=>X"00",
39537=>X"00",
39538=>X"00",
39539=>X"00",
39540=>X"00",
39541=>X"00",
39542=>X"00",
39543=>X"00",
39544=>X"00",
39545=>X"00",
39546=>X"00",
39547=>X"00",
39548=>X"00",
39549=>X"00",
39550=>X"00",
39551=>X"00",
39552=>X"00",
39553=>X"00",
39554=>X"00",
39555=>X"00",
39556=>X"00",
39557=>X"00",
39558=>X"00",
39559=>X"00",
39560=>X"00",
39561=>X"00",
39562=>X"00",
39563=>X"00",
39564=>X"00",
39565=>X"00",
39566=>X"00",
39567=>X"00",
39568=>X"00",
39569=>X"00",
39570=>X"00",
39571=>X"00",
39572=>X"00",
39573=>X"00",
39574=>X"00",
39575=>X"00",
39576=>X"00",
39577=>X"00",
39578=>X"00",
39579=>X"00",
39580=>X"00",
39581=>X"00",
39582=>X"00",
39583=>X"00",
39584=>X"00",
39585=>X"00",
39586=>X"00",
39587=>X"00",
39588=>X"00",
39589=>X"00",
39590=>X"00",
39591=>X"00",
39592=>X"00",
39593=>X"00",
39594=>X"00",
39595=>X"00",
39596=>X"00",
39597=>X"00",
39598=>X"00",
39599=>X"00",
39600=>X"00",
39601=>X"00",
39602=>X"00",
39603=>X"00",
39604=>X"00",
39605=>X"00",
39606=>X"00",
39607=>X"00",
39608=>X"00",
39609=>X"00",
39610=>X"00",
39611=>X"00",
39612=>X"00",
39613=>X"00",
39614=>X"00",
39615=>X"00",
39616=>X"00",
39617=>X"00",
39618=>X"00",
39619=>X"00",
39620=>X"00",
39621=>X"00",
39622=>X"00",
39623=>X"00",
39624=>X"00",
39625=>X"00",
39626=>X"00",
39627=>X"00",
39628=>X"00",
39629=>X"00",
39630=>X"00",
39631=>X"00",
39632=>X"00",
39633=>X"00",
39634=>X"00",
39635=>X"00",
39636=>X"00",
39637=>X"00",
39638=>X"00",
39639=>X"00",
39640=>X"00",
39641=>X"00",
39642=>X"00",
39643=>X"00",
39644=>X"00",
39645=>X"00",
39646=>X"00",
39647=>X"00",
39648=>X"00",
39649=>X"00",
39650=>X"00",
39651=>X"00",
39652=>X"00",
39653=>X"00",
39654=>X"00",
39655=>X"00",
39656=>X"00",
39657=>X"00",
39658=>X"00",
39659=>X"00",
39660=>X"00",
39661=>X"00",
39662=>X"00",
39663=>X"00",
39664=>X"00",
39665=>X"00",
39666=>X"00",
39667=>X"00",
39668=>X"00",
39669=>X"00",
39670=>X"00",
39671=>X"00",
39672=>X"00",
39673=>X"00",
39674=>X"00",
39675=>X"00",
39676=>X"00",
39677=>X"00",
39678=>X"00",
39679=>X"00",
39680=>X"00",
39681=>X"00",
39682=>X"00",
39683=>X"00",
39684=>X"00",
39685=>X"00",
39686=>X"00",
39687=>X"00",
39688=>X"00",
39689=>X"00",
39690=>X"00",
39691=>X"00",
39692=>X"00",
39693=>X"00",
39694=>X"00",
39695=>X"00",
39696=>X"00",
39697=>X"00",
39698=>X"00",
39699=>X"00",
39700=>X"00",
39701=>X"00",
39702=>X"00",
39703=>X"00",
39704=>X"00",
39705=>X"00",
39706=>X"00",
39707=>X"00",
39708=>X"00",
39709=>X"00",
39710=>X"00",
39711=>X"00",
39712=>X"00",
39713=>X"00",
39714=>X"00",
39715=>X"00",
39716=>X"00",
39717=>X"00",
39718=>X"00",
39719=>X"00",
39720=>X"00",
39721=>X"00",
39722=>X"00",
39723=>X"00",
39724=>X"00",
39725=>X"00",
39726=>X"00",
39727=>X"00",
39728=>X"00",
39729=>X"00",
39730=>X"00",
39731=>X"00",
39732=>X"00",
39733=>X"00",
39734=>X"00",
39735=>X"00",
39736=>X"00",
39737=>X"00",
39738=>X"00",
39739=>X"00",
39740=>X"00",
39741=>X"00",
39742=>X"00",
39743=>X"00",
39744=>X"00",
39745=>X"00",
39746=>X"00",
39747=>X"00",
39748=>X"00",
39749=>X"00",
39750=>X"00",
39751=>X"00",
39752=>X"00",
39753=>X"00",
39754=>X"00",
39755=>X"00",
39756=>X"00",
39757=>X"00",
39758=>X"00",
39759=>X"00",
39760=>X"00",
39761=>X"00",
39762=>X"00",
39763=>X"00",
39764=>X"00",
39765=>X"00",
39766=>X"00",
39767=>X"00",
39768=>X"00",
39769=>X"00",
39770=>X"00",
39771=>X"00",
39772=>X"00",
39773=>X"00",
39774=>X"00",
39775=>X"00",
39776=>X"00",
39777=>X"00",
39778=>X"00",
39779=>X"00",
39780=>X"00",
39781=>X"00",
39782=>X"00",
39783=>X"00",
39784=>X"00",
39785=>X"00",
39786=>X"00",
39787=>X"00",
39788=>X"00",
39789=>X"00",
39790=>X"00",
39791=>X"00",
39792=>X"00",
39793=>X"00",
39794=>X"00",
39795=>X"00",
39796=>X"00",
39797=>X"00",
39798=>X"00",
39799=>X"00",
39800=>X"00",
39801=>X"00",
39802=>X"00",
39803=>X"00",
39804=>X"00",
39805=>X"00",
39806=>X"00",
39807=>X"00",
39808=>X"00",
39809=>X"00",
39810=>X"00",
39811=>X"00",
39812=>X"00",
39813=>X"00",
39814=>X"00",
39815=>X"00",
39816=>X"00",
39817=>X"00",
39818=>X"00",
39819=>X"00",
39820=>X"00",
39821=>X"00",
39822=>X"00",
39823=>X"00",
39824=>X"00",
39825=>X"00",
39826=>X"00",
39827=>X"00",
39828=>X"00",
39829=>X"00",
39830=>X"00",
39831=>X"00",
39832=>X"00",
39833=>X"00",
39834=>X"00",
39835=>X"00",
39836=>X"00",
39837=>X"00",
39838=>X"00",
39839=>X"00",
39840=>X"00",
39841=>X"00",
39842=>X"00",
39843=>X"00",
39844=>X"00",
39845=>X"00",
39846=>X"00",
39847=>X"00",
39848=>X"00",
39849=>X"00",
39850=>X"00",
39851=>X"00",
39852=>X"00",
39853=>X"00",
39854=>X"00",
39855=>X"00",
39856=>X"00",
39857=>X"00",
39858=>X"00",
39859=>X"00",
39860=>X"00",
39861=>X"00",
39862=>X"00",
39863=>X"00",
39864=>X"00",
39865=>X"00",
39866=>X"00",
39867=>X"00",
39868=>X"00",
39869=>X"00",
39870=>X"00",
39871=>X"00",
39872=>X"00",
39873=>X"00",
39874=>X"00",
39875=>X"00",
39876=>X"00",
39877=>X"00",
39878=>X"00",
39879=>X"00",
39880=>X"00",
39881=>X"00",
39882=>X"00",
39883=>X"00",
39884=>X"00",
39885=>X"00",
39886=>X"00",
39887=>X"00",
39888=>X"00",
39889=>X"00",
39890=>X"00",
39891=>X"00",
39892=>X"00",
39893=>X"00",
39894=>X"00",
39895=>X"00",
39896=>X"00",
39897=>X"00",
39898=>X"00",
39899=>X"00",
39900=>X"00",
39901=>X"00",
39902=>X"00",
39903=>X"00",
39904=>X"00",
39905=>X"00",
39906=>X"00",
39907=>X"00",
39908=>X"00",
39909=>X"00",
39910=>X"00",
39911=>X"00",
39912=>X"00",
39913=>X"00",
39914=>X"00",
39915=>X"00",
39916=>X"00",
39917=>X"00",
39918=>X"00",
39919=>X"00",
39920=>X"00",
39921=>X"00",
39922=>X"00",
39923=>X"00",
39924=>X"00",
39925=>X"00",
39926=>X"00",
39927=>X"00",
39928=>X"00",
39929=>X"00",
39930=>X"00",
39931=>X"00",
39932=>X"00",
39933=>X"00",
39934=>X"00",
39935=>X"00",
39936=>X"00",
39937=>X"00",
39938=>X"00",
39939=>X"00",
39940=>X"00",
39941=>X"00",
39942=>X"00",
39943=>X"00",
39944=>X"00",
39945=>X"00",
39946=>X"00",
39947=>X"00",
39948=>X"00",
39949=>X"00",
39950=>X"00",
39951=>X"00",
39952=>X"00",
39953=>X"00",
39954=>X"00",
39955=>X"00",
39956=>X"00",
39957=>X"00",
39958=>X"00",
39959=>X"00",
39960=>X"00",
39961=>X"00",
39962=>X"00",
39963=>X"00",
39964=>X"00",
39965=>X"00",
39966=>X"00",
39967=>X"00",
39968=>X"00",
39969=>X"00",
39970=>X"00",
39971=>X"00",
39972=>X"00",
39973=>X"00",
39974=>X"00",
39975=>X"00",
39976=>X"00",
39977=>X"00",
39978=>X"00",
39979=>X"00",
39980=>X"00",
39981=>X"00",
39982=>X"00",
39983=>X"00",
39984=>X"00",
39985=>X"00",
39986=>X"00",
39987=>X"00",
39988=>X"00",
39989=>X"00",
39990=>X"00",
39991=>X"00",
39992=>X"00",
39993=>X"00",
39994=>X"00",
39995=>X"00",
39996=>X"00",
39997=>X"00",
39998=>X"00",
39999=>X"00",
40000=>X"00",
40001=>X"00",
40002=>X"00",
40003=>X"00",
40004=>X"00",
40005=>X"00",
40006=>X"00",
40007=>X"00",
40008=>X"00",
40009=>X"00",
40010=>X"00",
40011=>X"00",
40012=>X"00",
40013=>X"00",
40014=>X"00",
40015=>X"00",
40016=>X"00",
40017=>X"00",
40018=>X"00",
40019=>X"00",
40020=>X"00",
40021=>X"00",
40022=>X"00",
40023=>X"00",
40024=>X"00",
40025=>X"00",
40026=>X"00",
40027=>X"00",
40028=>X"00",
40029=>X"00",
40030=>X"00",
40031=>X"00",
40032=>X"00",
40033=>X"00",
40034=>X"00",
40035=>X"00",
40036=>X"00",
40037=>X"00",
40038=>X"00",
40039=>X"00",
40040=>X"00",
40041=>X"00",
40042=>X"00",
40043=>X"00",
40044=>X"00",
40045=>X"00",
40046=>X"00",
40047=>X"00",
40048=>X"00",
40049=>X"00",
40050=>X"00",
40051=>X"00",
40052=>X"00",
40053=>X"00",
40054=>X"00",
40055=>X"00",
40056=>X"00",
40057=>X"00",
40058=>X"00",
40059=>X"00",
40060=>X"00",
40061=>X"00",
40062=>X"00",
40063=>X"00",
40064=>X"00",
40065=>X"00",
40066=>X"00",
40067=>X"00",
40068=>X"00",
40069=>X"00",
40070=>X"00",
40071=>X"00",
40072=>X"00",
40073=>X"00",
40074=>X"00",
40075=>X"00",
40076=>X"00",
40077=>X"00",
40078=>X"00",
40079=>X"00",
40080=>X"00",
40081=>X"00",
40082=>X"00",
40083=>X"00",
40084=>X"00",
40085=>X"00",
40086=>X"00",
40087=>X"00",
40088=>X"00",
40089=>X"00",
40090=>X"00",
40091=>X"00",
40092=>X"00",
40093=>X"00",
40094=>X"00",
40095=>X"00",
40096=>X"00",
40097=>X"00",
40098=>X"00",
40099=>X"00",
40100=>X"00",
40101=>X"00",
40102=>X"00",
40103=>X"00",
40104=>X"00",
40105=>X"00",
40106=>X"00",
40107=>X"00",
40108=>X"00",
40109=>X"00",
40110=>X"00",
40111=>X"00",
40112=>X"00",
40113=>X"00",
40114=>X"00",
40115=>X"00",
40116=>X"00",
40117=>X"00",
40118=>X"00",
40119=>X"00",
40120=>X"00",
40121=>X"00",
40122=>X"00",
40123=>X"00",
40124=>X"00",
40125=>X"00",
40126=>X"00",
40127=>X"00",
40128=>X"00",
40129=>X"00",
40130=>X"00",
40131=>X"00",
40132=>X"00",
40133=>X"00",
40134=>X"00",
40135=>X"00",
40136=>X"00",
40137=>X"00",
40138=>X"00",
40139=>X"00",
40140=>X"00",
40141=>X"00",
40142=>X"00",
40143=>X"00",
40144=>X"00",
40145=>X"00",
40146=>X"00",
40147=>X"00",
40148=>X"00",
40149=>X"00",
40150=>X"00",
40151=>X"00",
40152=>X"00",
40153=>X"00",
40154=>X"00",
40155=>X"00",
40156=>X"00",
40157=>X"00",
40158=>X"00",
40159=>X"00",
40160=>X"00",
40161=>X"00",
40162=>X"00",
40163=>X"00",
40164=>X"00",
40165=>X"00",
40166=>X"00",
40167=>X"00",
40168=>X"00",
40169=>X"00",
40170=>X"00",
40171=>X"00",
40172=>X"00",
40173=>X"00",
40174=>X"00",
40175=>X"00",
40176=>X"00",
40177=>X"00",
40178=>X"00",
40179=>X"00",
40180=>X"00",
40181=>X"00",
40182=>X"00",
40183=>X"00",
40184=>X"00",
40185=>X"00",
40186=>X"00",
40187=>X"00",
40188=>X"00",
40189=>X"00",
40190=>X"00",
40191=>X"00",
40192=>X"00",
40193=>X"00",
40194=>X"00",
40195=>X"00",
40196=>X"00",
40197=>X"00",
40198=>X"00",
40199=>X"00",
40200=>X"00",
40201=>X"00",
40202=>X"00",
40203=>X"00",
40204=>X"00",
40205=>X"00",
40206=>X"00",
40207=>X"00",
40208=>X"00",
40209=>X"00",
40210=>X"00",
40211=>X"00",
40212=>X"00",
40213=>X"00",
40214=>X"00",
40215=>X"00",
40216=>X"00",
40217=>X"00",
40218=>X"00",
40219=>X"00",
40220=>X"00",
40221=>X"00",
40222=>X"00",
40223=>X"00",
40224=>X"00",
40225=>X"00",
40226=>X"00",
40227=>X"00",
40228=>X"00",
40229=>X"00",
40230=>X"00",
40231=>X"00",
40232=>X"00",
40233=>X"00",
40234=>X"00",
40235=>X"00",
40236=>X"00",
40237=>X"00",
40238=>X"00",
40239=>X"00",
40240=>X"00",
40241=>X"00",
40242=>X"00",
40243=>X"00",
40244=>X"00",
40245=>X"00",
40246=>X"00",
40247=>X"00",
40248=>X"00",
40249=>X"00",
40250=>X"00",
40251=>X"00",
40252=>X"00",
40253=>X"00",
40254=>X"00",
40255=>X"00",
40256=>X"00",
40257=>X"00",
40258=>X"00",
40259=>X"00",
40260=>X"00",
40261=>X"00",
40262=>X"00",
40263=>X"00",
40264=>X"00",
40265=>X"00",
40266=>X"00",
40267=>X"00",
40268=>X"00",
40269=>X"00",
40270=>X"00",
40271=>X"00",
40272=>X"00",
40273=>X"00",
40274=>X"00",
40275=>X"00",
40276=>X"00",
40277=>X"00",
40278=>X"00",
40279=>X"00",
40280=>X"00",
40281=>X"00",
40282=>X"00",
40283=>X"00",
40284=>X"00",
40285=>X"00",
40286=>X"00",
40287=>X"00",
40288=>X"00",
40289=>X"00",
40290=>X"00",
40291=>X"00",
40292=>X"00",
40293=>X"00",
40294=>X"00",
40295=>X"00",
40296=>X"00",
40297=>X"00",
40298=>X"00",
40299=>X"00",
40300=>X"00",
40301=>X"00",
40302=>X"00",
40303=>X"00",
40304=>X"00",
40305=>X"00",
40306=>X"00",
40307=>X"00",
40308=>X"00",
40309=>X"00",
40310=>X"00",
40311=>X"00",
40312=>X"00",
40313=>X"00",
40314=>X"00",
40315=>X"00",
40316=>X"00",
40317=>X"00",
40318=>X"00",
40319=>X"00",
40320=>X"00",
40321=>X"00",
40322=>X"00",
40323=>X"00",
40324=>X"00",
40325=>X"00",
40326=>X"00",
40327=>X"00",
40328=>X"00",
40329=>X"00",
40330=>X"00",
40331=>X"00",
40332=>X"00",
40333=>X"00",
40334=>X"00",
40335=>X"00",
40336=>X"00",
40337=>X"00",
40338=>X"00",
40339=>X"00",
40340=>X"00",
40341=>X"00",
40342=>X"00",
40343=>X"00",
40344=>X"00",
40345=>X"00",
40346=>X"00",
40347=>X"00",
40348=>X"00",
40349=>X"00",
40350=>X"00",
40351=>X"00",
40352=>X"00",
40353=>X"00",
40354=>X"00",
40355=>X"00",
40356=>X"00",
40357=>X"00",
40358=>X"00",
40359=>X"00",
40360=>X"00",
40361=>X"00",
40362=>X"00",
40363=>X"00",
40364=>X"00",
40365=>X"00",
40366=>X"00",
40367=>X"00",
40368=>X"00",
40369=>X"00",
40370=>X"00",
40371=>X"00",
40372=>X"00",
40373=>X"00",
40374=>X"00",
40375=>X"00",
40376=>X"00",
40377=>X"00",
40378=>X"00",
40379=>X"00",
40380=>X"00",
40381=>X"00",
40382=>X"00",
40383=>X"00",
40384=>X"00",
40385=>X"00",
40386=>X"00",
40387=>X"00",
40388=>X"00",
40389=>X"00",
40390=>X"00",
40391=>X"00",
40392=>X"00",
40393=>X"00",
40394=>X"00",
40395=>X"00",
40396=>X"00",
40397=>X"00",
40398=>X"00",
40399=>X"00",
40400=>X"00",
40401=>X"00",
40402=>X"00",
40403=>X"00",
40404=>X"00",
40405=>X"00",
40406=>X"00",
40407=>X"00",
40408=>X"00",
40409=>X"00",
40410=>X"00",
40411=>X"00",
40412=>X"00",
40413=>X"00",
40414=>X"00",
40415=>X"00",
40416=>X"00",
40417=>X"00",
40418=>X"00",
40419=>X"00",
40420=>X"00",
40421=>X"00",
40422=>X"00",
40423=>X"00",
40424=>X"00",
40425=>X"00",
40426=>X"00",
40427=>X"00",
40428=>X"00",
40429=>X"00",
40430=>X"00",
40431=>X"00",
40432=>X"00",
40433=>X"00",
40434=>X"00",
40435=>X"00",
40436=>X"00",
40437=>X"00",
40438=>X"00",
40439=>X"00",
40440=>X"00",
40441=>X"00",
40442=>X"00",
40443=>X"00",
40444=>X"00",
40445=>X"00",
40446=>X"00",
40447=>X"00",
40448=>X"00",
40449=>X"00",
40450=>X"00",
40451=>X"00",
40452=>X"00",
40453=>X"00",
40454=>X"00",
40455=>X"00",
40456=>X"00",
40457=>X"00",
40458=>X"00",
40459=>X"00",
40460=>X"00",
40461=>X"00",
40462=>X"00",
40463=>X"00",
40464=>X"00",
40465=>X"00",
40466=>X"00",
40467=>X"00",
40468=>X"00",
40469=>X"00",
40470=>X"00",
40471=>X"00",
40472=>X"00",
40473=>X"00",
40474=>X"00",
40475=>X"00",
40476=>X"00",
40477=>X"00",
40478=>X"00",
40479=>X"00",
40480=>X"00",
40481=>X"00",
40482=>X"00",
40483=>X"00",
40484=>X"00",
40485=>X"00",
40486=>X"00",
40487=>X"00",
40488=>X"00",
40489=>X"00",
40490=>X"00",
40491=>X"00",
40492=>X"00",
40493=>X"00",
40494=>X"00",
40495=>X"00",
40496=>X"00",
40497=>X"00",
40498=>X"00",
40499=>X"00",
40500=>X"00",
40501=>X"00",
40502=>X"00",
40503=>X"00",
40504=>X"00",
40505=>X"00",
40506=>X"00",
40507=>X"00",
40508=>X"00",
40509=>X"00",
40510=>X"00",
40511=>X"00",
40512=>X"00",
40513=>X"00",
40514=>X"00",
40515=>X"00",
40516=>X"00",
40517=>X"00",
40518=>X"00",
40519=>X"00",
40520=>X"00",
40521=>X"00",
40522=>X"00",
40523=>X"00",
40524=>X"00",
40525=>X"00",
40526=>X"00",
40527=>X"00",
40528=>X"00",
40529=>X"00",
40530=>X"00",
40531=>X"00",
40532=>X"00",
40533=>X"00",
40534=>X"00",
40535=>X"00",
40536=>X"00",
40537=>X"00",
40538=>X"00",
40539=>X"00",
40540=>X"00",
40541=>X"00",
40542=>X"00",
40543=>X"00",
40544=>X"00",
40545=>X"00",
40546=>X"00",
40547=>X"00",
40548=>X"00",
40549=>X"00",
40550=>X"00",
40551=>X"00",
40552=>X"00",
40553=>X"00",
40554=>X"00",
40555=>X"00",
40556=>X"00",
40557=>X"00",
40558=>X"00",
40559=>X"00",
40560=>X"00",
40561=>X"00",
40562=>X"00",
40563=>X"00",
40564=>X"00",
40565=>X"00",
40566=>X"00",
40567=>X"00",
40568=>X"00",
40569=>X"00",
40570=>X"00",
40571=>X"00",
40572=>X"00",
40573=>X"00",
40574=>X"00",
40575=>X"00",
40576=>X"00",
40577=>X"00",
40578=>X"00",
40579=>X"00",
40580=>X"00",
40581=>X"00",
40582=>X"00",
40583=>X"00",
40584=>X"00",
40585=>X"00",
40586=>X"00",
40587=>X"00",
40588=>X"00",
40589=>X"00",
40590=>X"00",
40591=>X"00",
40592=>X"00",
40593=>X"00",
40594=>X"00",
40595=>X"00",
40596=>X"00",
40597=>X"00",
40598=>X"00",
40599=>X"00",
40600=>X"00",
40601=>X"00",
40602=>X"00",
40603=>X"00",
40604=>X"00",
40605=>X"00",
40606=>X"00",
40607=>X"00",
40608=>X"00",
40609=>X"00",
40610=>X"00",
40611=>X"00",
40612=>X"00",
40613=>X"00",
40614=>X"00",
40615=>X"00",
40616=>X"00",
40617=>X"00",
40618=>X"00",
40619=>X"00",
40620=>X"00",
40621=>X"00",
40622=>X"00",
40623=>X"00",
40624=>X"00",
40625=>X"00",
40626=>X"00",
40627=>X"00",
40628=>X"00",
40629=>X"00",
40630=>X"00",
40631=>X"00",
40632=>X"00",
40633=>X"00",
40634=>X"00",
40635=>X"00",
40636=>X"00",
40637=>X"00",
40638=>X"00",
40639=>X"00",
40640=>X"00",
40641=>X"00",
40642=>X"00",
40643=>X"00",
40644=>X"00",
40645=>X"00",
40646=>X"00",
40647=>X"00",
40648=>X"00",
40649=>X"00",
40650=>X"00",
40651=>X"00",
40652=>X"00",
40653=>X"00",
40654=>X"00",
40655=>X"00",
40656=>X"00",
40657=>X"00",
40658=>X"00",
40659=>X"00",
40660=>X"00",
40661=>X"00",
40662=>X"00",
40663=>X"00",
40664=>X"00",
40665=>X"00",
40666=>X"00",
40667=>X"00",
40668=>X"00",
40669=>X"00",
40670=>X"00",
40671=>X"00",
40672=>X"00",
40673=>X"00",
40674=>X"00",
40675=>X"00",
40676=>X"00",
40677=>X"00",
40678=>X"00",
40679=>X"00",
40680=>X"00",
40681=>X"00",
40682=>X"00",
40683=>X"00",
40684=>X"00",
40685=>X"00",
40686=>X"00",
40687=>X"00",
40688=>X"00",
40689=>X"00",
40690=>X"00",
40691=>X"00",
40692=>X"00",
40693=>X"00",
40694=>X"00",
40695=>X"00",
40696=>X"00",
40697=>X"00",
40698=>X"00",
40699=>X"00",
40700=>X"00",
40701=>X"00",
40702=>X"00",
40703=>X"00",
40704=>X"00",
40705=>X"00",
40706=>X"00",
40707=>X"00",
40708=>X"00",
40709=>X"00",
40710=>X"00",
40711=>X"00",
40712=>X"00",
40713=>X"00",
40714=>X"00",
40715=>X"00",
40716=>X"00",
40717=>X"00",
40718=>X"00",
40719=>X"00",
40720=>X"00",
40721=>X"00",
40722=>X"00",
40723=>X"00",
40724=>X"00",
40725=>X"00",
40726=>X"00",
40727=>X"00",
40728=>X"00",
40729=>X"00",
40730=>X"00",
40731=>X"00",
40732=>X"00",
40733=>X"00",
40734=>X"00",
40735=>X"00",
40736=>X"00",
40737=>X"00",
40738=>X"00",
40739=>X"00",
40740=>X"00",
40741=>X"00",
40742=>X"00",
40743=>X"00",
40744=>X"00",
40745=>X"00",
40746=>X"00",
40747=>X"00",
40748=>X"00",
40749=>X"00",
40750=>X"00",
40751=>X"00",
40752=>X"00",
40753=>X"00",
40754=>X"00",
40755=>X"00",
40756=>X"00",
40757=>X"00",
40758=>X"00",
40759=>X"00",
40760=>X"00",
40761=>X"00",
40762=>X"00",
40763=>X"00",
40764=>X"00",
40765=>X"00",
40766=>X"00",
40767=>X"00",
40768=>X"00",
40769=>X"00",
40770=>X"00",
40771=>X"00",
40772=>X"00",
40773=>X"00",
40774=>X"00",
40775=>X"00",
40776=>X"00",
40777=>X"00",
40778=>X"00",
40779=>X"00",
40780=>X"00",
40781=>X"00",
40782=>X"00",
40783=>X"00",
40784=>X"00",
40785=>X"00",
40786=>X"00",
40787=>X"00",
40788=>X"00",
40789=>X"00",
40790=>X"00",
40791=>X"00",
40792=>X"00",
40793=>X"00",
40794=>X"00",
40795=>X"00",
40796=>X"00",
40797=>X"00",
40798=>X"00",
40799=>X"00",
40800=>X"00",
40801=>X"00",
40802=>X"00",
40803=>X"00",
40804=>X"00",
40805=>X"00",
40806=>X"00",
40807=>X"00",
40808=>X"00",
40809=>X"00",
40810=>X"00",
40811=>X"00",
40812=>X"00",
40813=>X"00",
40814=>X"00",
40815=>X"00",
40816=>X"00",
40817=>X"00",
40818=>X"00",
40819=>X"00",
40820=>X"00",
40821=>X"00",
40822=>X"00",
40823=>X"00",
40824=>X"00",
40825=>X"00",
40826=>X"00",
40827=>X"00",
40828=>X"00",
40829=>X"00",
40830=>X"00",
40831=>X"00",
40832=>X"00",
40833=>X"00",
40834=>X"00",
40835=>X"00",
40836=>X"00",
40837=>X"00",
40838=>X"00",
40839=>X"00",
40840=>X"00",
40841=>X"00",
40842=>X"00",
40843=>X"00",
40844=>X"00",
40845=>X"00",
40846=>X"00",
40847=>X"00",
40848=>X"00",
40849=>X"00",
40850=>X"00",
40851=>X"00",
40852=>X"00",
40853=>X"00",
40854=>X"00",
40855=>X"00",
40856=>X"00",
40857=>X"00",
40858=>X"00",
40859=>X"00",
40860=>X"00",
40861=>X"00",
40862=>X"00",
40863=>X"00",
40864=>X"00",
40865=>X"00",
40866=>X"00",
40867=>X"00",
40868=>X"00",
40869=>X"00",
40870=>X"00",
40871=>X"00",
40872=>X"00",
40873=>X"00",
40874=>X"00",
40875=>X"00",
40876=>X"00",
40877=>X"00",
40878=>X"00",
40879=>X"00",
40880=>X"00",
40881=>X"00",
40882=>X"00",
40883=>X"00",
40884=>X"00",
40885=>X"00",
40886=>X"00",
40887=>X"00",
40888=>X"00",
40889=>X"00",
40890=>X"00",
40891=>X"00",
40892=>X"00",
40893=>X"00",
40894=>X"00",
40895=>X"00",
40896=>X"00",
40897=>X"00",
40898=>X"00",
40899=>X"00",
40900=>X"00",
40901=>X"00",
40902=>X"00",
40903=>X"00",
40904=>X"00",
40905=>X"00",
40906=>X"00",
40907=>X"00",
40908=>X"00",
40909=>X"00",
40910=>X"00",
40911=>X"00",
40912=>X"00",
40913=>X"00",
40914=>X"00",
40915=>X"00",
40916=>X"00",
40917=>X"00",
40918=>X"00",
40919=>X"00",
40920=>X"00",
40921=>X"00",
40922=>X"00",
40923=>X"00",
40924=>X"00",
40925=>X"00",
40926=>X"00",
40927=>X"00",
40928=>X"00",
40929=>X"00",
40930=>X"00",
40931=>X"00",
40932=>X"00",
40933=>X"00",
40934=>X"00",
40935=>X"00",
40936=>X"00",
40937=>X"00",
40938=>X"00",
40939=>X"00",
40940=>X"00",
40941=>X"00",
40942=>X"00",
40943=>X"00",
40944=>X"00",
40945=>X"00",
40946=>X"00",
40947=>X"00",
40948=>X"00",
40949=>X"00",
40950=>X"00",
40951=>X"00",
40952=>X"00",
40953=>X"00",
40954=>X"00",
40955=>X"00",
40956=>X"00",
40957=>X"00",
40958=>X"00",
40959=>X"00",
40960=>X"00",
40961=>X"00",
40962=>X"00",
40963=>X"00",
40964=>X"00",
40965=>X"00",
40966=>X"00",
40967=>X"00",
40968=>X"00",
40969=>X"00",
40970=>X"00",
40971=>X"00",
40972=>X"00",
40973=>X"00",
40974=>X"00",
40975=>X"00",
40976=>X"00",
40977=>X"00",
40978=>X"00",
40979=>X"00",
40980=>X"00",
40981=>X"00",
40982=>X"00",
40983=>X"00",
40984=>X"00",
40985=>X"00",
40986=>X"00",
40987=>X"00",
40988=>X"00",
40989=>X"00",
40990=>X"00",
40991=>X"00",
40992=>X"00",
40993=>X"00",
40994=>X"00",
40995=>X"00",
40996=>X"00",
40997=>X"00",
40998=>X"00",
40999=>X"00",
41000=>X"00",
41001=>X"00",
41002=>X"00",
41003=>X"00",
41004=>X"00",
41005=>X"00",
41006=>X"00",
41007=>X"00",
41008=>X"00",
41009=>X"00",
41010=>X"00",
41011=>X"00",
41012=>X"00",
41013=>X"00",
41014=>X"00",
41015=>X"00",
41016=>X"00",
41017=>X"00",
41018=>X"00",
41019=>X"00",
41020=>X"00",
41021=>X"00",
41022=>X"00",
41023=>X"00",
41024=>X"00",
41025=>X"00",
41026=>X"00",
41027=>X"00",
41028=>X"00",
41029=>X"00",
41030=>X"00",
41031=>X"00",
41032=>X"00",
41033=>X"00",
41034=>X"00",
41035=>X"00",
41036=>X"00",
41037=>X"00",
41038=>X"00",
41039=>X"00",
41040=>X"00",
41041=>X"00",
41042=>X"00",
41043=>X"00",
41044=>X"00",
41045=>X"00",
41046=>X"00",
41047=>X"00",
41048=>X"00",
41049=>X"00",
41050=>X"00",
41051=>X"00",
41052=>X"00",
41053=>X"00",
41054=>X"00",
41055=>X"00",
41056=>X"00",
41057=>X"00",
41058=>X"00",
41059=>X"00",
41060=>X"00",
41061=>X"00",
41062=>X"00",
41063=>X"00",
41064=>X"00",
41065=>X"00",
41066=>X"00",
41067=>X"00",
41068=>X"00",
41069=>X"00",
41070=>X"00",
41071=>X"00",
41072=>X"00",
41073=>X"00",
41074=>X"00",
41075=>X"00",
41076=>X"00",
41077=>X"00",
41078=>X"00",
41079=>X"00",
41080=>X"00",
41081=>X"00",
41082=>X"00",
41083=>X"00",
41084=>X"00",
41085=>X"00",
41086=>X"00",
41087=>X"00",
41088=>X"00",
41089=>X"00",
41090=>X"00",
41091=>X"00",
41092=>X"00",
41093=>X"00",
41094=>X"00",
41095=>X"00",
41096=>X"00",
41097=>X"00",
41098=>X"00",
41099=>X"00",
41100=>X"00",
41101=>X"00",
41102=>X"00",
41103=>X"00",
41104=>X"00",
41105=>X"00",
41106=>X"00",
41107=>X"00",
41108=>X"00",
41109=>X"00",
41110=>X"00",
41111=>X"00",
41112=>X"00",
41113=>X"00",
41114=>X"00",
41115=>X"00",
41116=>X"00",
41117=>X"00",
41118=>X"00",
41119=>X"00",
41120=>X"00",
41121=>X"00",
41122=>X"00",
41123=>X"00",
41124=>X"00",
41125=>X"00",
41126=>X"00",
41127=>X"00",
41128=>X"00",
41129=>X"00",
41130=>X"00",
41131=>X"00",
41132=>X"00",
41133=>X"00",
41134=>X"00",
41135=>X"00",
41136=>X"00",
41137=>X"00",
41138=>X"00",
41139=>X"00",
41140=>X"00",
41141=>X"00",
41142=>X"00",
41143=>X"00",
41144=>X"00",
41145=>X"00",
41146=>X"00",
41147=>X"00",
41148=>X"00",
41149=>X"00",
41150=>X"00",
41151=>X"00",
41152=>X"00",
41153=>X"00",
41154=>X"00",
41155=>X"00",
41156=>X"00",
41157=>X"00",
41158=>X"00",
41159=>X"00",
41160=>X"00",
41161=>X"00",
41162=>X"00",
41163=>X"00",
41164=>X"00",
41165=>X"00",
41166=>X"00",
41167=>X"00",
41168=>X"00",
41169=>X"00",
41170=>X"00",
41171=>X"00",
41172=>X"00",
41173=>X"00",
41174=>X"00",
41175=>X"00",
41176=>X"00",
41177=>X"00",
41178=>X"00",
41179=>X"00",
41180=>X"00",
41181=>X"00",
41182=>X"00",
41183=>X"00",
41184=>X"00",
41185=>X"00",
41186=>X"00",
41187=>X"00",
41188=>X"00",
41189=>X"00",
41190=>X"00",
41191=>X"00",
41192=>X"00",
41193=>X"00",
41194=>X"00",
41195=>X"00",
41196=>X"00",
41197=>X"00",
41198=>X"00",
41199=>X"00",
41200=>X"00",
41201=>X"00",
41202=>X"00",
41203=>X"00",
41204=>X"00",
41205=>X"00",
41206=>X"00",
41207=>X"00",
41208=>X"00",
41209=>X"00",
41210=>X"00",
41211=>X"00",
41212=>X"00",
41213=>X"00",
41214=>X"00",
41215=>X"00",
41216=>X"00",
41217=>X"00",
41218=>X"00",
41219=>X"00",
41220=>X"00",
41221=>X"00",
41222=>X"00",
41223=>X"00",
41224=>X"00",
41225=>X"00",
41226=>X"00",
41227=>X"00",
41228=>X"00",
41229=>X"00",
41230=>X"00",
41231=>X"00",
41232=>X"00",
41233=>X"00",
41234=>X"00",
41235=>X"00",
41236=>X"00",
41237=>X"00",
41238=>X"00",
41239=>X"00",
41240=>X"00",
41241=>X"00",
41242=>X"00",
41243=>X"00",
41244=>X"00",
41245=>X"00",
41246=>X"00",
41247=>X"00",
41248=>X"00",
41249=>X"00",
41250=>X"00",
41251=>X"00",
41252=>X"00",
41253=>X"00",
41254=>X"00",
41255=>X"00",
41256=>X"00",
41257=>X"00",
41258=>X"00",
41259=>X"00",
41260=>X"00",
41261=>X"00",
41262=>X"00",
41263=>X"00",
41264=>X"00",
41265=>X"00",
41266=>X"00",
41267=>X"00",
41268=>X"00",
41269=>X"00",
41270=>X"00",
41271=>X"00",
41272=>X"00",
41273=>X"00",
41274=>X"00",
41275=>X"00",
41276=>X"00",
41277=>X"00",
41278=>X"00",
41279=>X"00",
41280=>X"00",
41281=>X"00",
41282=>X"00",
41283=>X"00",
41284=>X"00",
41285=>X"00",
41286=>X"00",
41287=>X"00",
41288=>X"00",
41289=>X"00",
41290=>X"00",
41291=>X"00",
41292=>X"00",
41293=>X"00",
41294=>X"00",
41295=>X"00",
41296=>X"00",
41297=>X"00",
41298=>X"00",
41299=>X"00",
41300=>X"00",
41301=>X"00",
41302=>X"00",
41303=>X"00",
41304=>X"00",
41305=>X"00",
41306=>X"00",
41307=>X"00",
41308=>X"00",
41309=>X"00",
41310=>X"00",
41311=>X"00",
41312=>X"00",
41313=>X"00",
41314=>X"00",
41315=>X"00",
41316=>X"00",
41317=>X"00",
41318=>X"00",
41319=>X"00",
41320=>X"00",
41321=>X"00",
41322=>X"00",
41323=>X"00",
41324=>X"00",
41325=>X"00",
41326=>X"00",
41327=>X"00",
41328=>X"00",
41329=>X"00",
41330=>X"00",
41331=>X"00",
41332=>X"00",
41333=>X"00",
41334=>X"00",
41335=>X"00",
41336=>X"00",
41337=>X"00",
41338=>X"00",
41339=>X"00",
41340=>X"00",
41341=>X"00",
41342=>X"00",
41343=>X"00",
41344=>X"00",
41345=>X"00",
41346=>X"00",
41347=>X"00",
41348=>X"00",
41349=>X"00",
41350=>X"00",
41351=>X"00",
41352=>X"00",
41353=>X"00",
41354=>X"00",
41355=>X"00",
41356=>X"00",
41357=>X"00",
41358=>X"00",
41359=>X"00",
41360=>X"00",
41361=>X"00",
41362=>X"00",
41363=>X"00",
41364=>X"00",
41365=>X"00",
41366=>X"00",
41367=>X"00",
41368=>X"00",
41369=>X"00",
41370=>X"00",
41371=>X"00",
41372=>X"00",
41373=>X"00",
41374=>X"00",
41375=>X"00",
41376=>X"00",
41377=>X"00",
41378=>X"00",
41379=>X"00",
41380=>X"00",
41381=>X"00",
41382=>X"00",
41383=>X"00",
41384=>X"00",
41385=>X"00",
41386=>X"00",
41387=>X"00",
41388=>X"00",
41389=>X"00",
41390=>X"00",
41391=>X"00",
41392=>X"00",
41393=>X"00",
41394=>X"00",
41395=>X"00",
41396=>X"00",
41397=>X"00",
41398=>X"00",
41399=>X"00",
41400=>X"00",
41401=>X"00",
41402=>X"00",
41403=>X"00",
41404=>X"00",
41405=>X"00",
41406=>X"00",
41407=>X"00",
41408=>X"00",
41409=>X"00",
41410=>X"00",
41411=>X"00",
41412=>X"00",
41413=>X"00",
41414=>X"00",
41415=>X"00",
41416=>X"00",
41417=>X"00",
41418=>X"00",
41419=>X"00",
41420=>X"00",
41421=>X"00",
41422=>X"00",
41423=>X"00",
41424=>X"00",
41425=>X"00",
41426=>X"00",
41427=>X"00",
41428=>X"00",
41429=>X"00",
41430=>X"00",
41431=>X"00",
41432=>X"00",
41433=>X"00",
41434=>X"00",
41435=>X"00",
41436=>X"00",
41437=>X"00",
41438=>X"00",
41439=>X"00",
41440=>X"00",
41441=>X"00",
41442=>X"00",
41443=>X"00",
41444=>X"00",
41445=>X"00",
41446=>X"00",
41447=>X"00",
41448=>X"00",
41449=>X"00",
41450=>X"00",
41451=>X"00",
41452=>X"00",
41453=>X"00",
41454=>X"00",
41455=>X"00",
41456=>X"00",
41457=>X"00",
41458=>X"00",
41459=>X"00",
41460=>X"00",
41461=>X"00",
41462=>X"00",
41463=>X"00",
41464=>X"00",
41465=>X"00",
41466=>X"00",
41467=>X"00",
41468=>X"00",
41469=>X"00",
41470=>X"00",
41471=>X"00",
41472=>X"00",
41473=>X"00",
41474=>X"00",
41475=>X"00",
41476=>X"00",
41477=>X"00",
41478=>X"00",
41479=>X"00",
41480=>X"00",
41481=>X"00",
41482=>X"00",
41483=>X"00",
41484=>X"00",
41485=>X"00",
41486=>X"00",
41487=>X"00",
41488=>X"00",
41489=>X"00",
41490=>X"00",
41491=>X"00",
41492=>X"00",
41493=>X"00",
41494=>X"00",
41495=>X"00",
41496=>X"00",
41497=>X"00",
41498=>X"00",
41499=>X"00",
41500=>X"00",
41501=>X"00",
41502=>X"00",
41503=>X"00",
41504=>X"00",
41505=>X"00",
41506=>X"00",
41507=>X"00",
41508=>X"00",
41509=>X"00",
41510=>X"00",
41511=>X"00",
41512=>X"00",
41513=>X"00",
41514=>X"00",
41515=>X"00",
41516=>X"00",
41517=>X"00",
41518=>X"00",
41519=>X"00",
41520=>X"00",
41521=>X"00",
41522=>X"00",
41523=>X"00",
41524=>X"00",
41525=>X"00",
41526=>X"00",
41527=>X"00",
41528=>X"00",
41529=>X"00",
41530=>X"00",
41531=>X"00",
41532=>X"00",
41533=>X"00",
41534=>X"00",
41535=>X"00",
41536=>X"00",
41537=>X"00",
41538=>X"00",
41539=>X"00",
41540=>X"00",
41541=>X"00",
41542=>X"00",
41543=>X"00",
41544=>X"00",
41545=>X"00",
41546=>X"00",
41547=>X"00",
41548=>X"00",
41549=>X"00",
41550=>X"00",
41551=>X"00",
41552=>X"00",
41553=>X"00",
41554=>X"00",
41555=>X"00",
41556=>X"00",
41557=>X"00",
41558=>X"00",
41559=>X"00",
41560=>X"00",
41561=>X"00",
41562=>X"00",
41563=>X"00",
41564=>X"00",
41565=>X"00",
41566=>X"00",
41567=>X"00",
41568=>X"00",
41569=>X"00",
41570=>X"00",
41571=>X"00",
41572=>X"00",
41573=>X"00",
41574=>X"00",
41575=>X"00",
41576=>X"00",
41577=>X"00",
41578=>X"00",
41579=>X"00",
41580=>X"00",
41581=>X"00",
41582=>X"00",
41583=>X"00",
41584=>X"00",
41585=>X"00",
41586=>X"00",
41587=>X"00",
41588=>X"00",
41589=>X"00",
41590=>X"00",
41591=>X"00",
41592=>X"00",
41593=>X"00",
41594=>X"00",
41595=>X"00",
41596=>X"00",
41597=>X"00",
41598=>X"00",
41599=>X"00",
41600=>X"00",
41601=>X"00",
41602=>X"00",
41603=>X"00",
41604=>X"00",
41605=>X"00",
41606=>X"00",
41607=>X"00",
41608=>X"00",
41609=>X"00",
41610=>X"00",
41611=>X"00",
41612=>X"00",
41613=>X"00",
41614=>X"00",
41615=>X"00",
41616=>X"00",
41617=>X"00",
41618=>X"00",
41619=>X"00",
41620=>X"00",
41621=>X"00",
41622=>X"00",
41623=>X"00",
41624=>X"00",
41625=>X"00",
41626=>X"00",
41627=>X"00",
41628=>X"00",
41629=>X"00",
41630=>X"00",
41631=>X"00",
41632=>X"00",
41633=>X"00",
41634=>X"00",
41635=>X"00",
41636=>X"00",
41637=>X"00",
41638=>X"00",
41639=>X"00",
41640=>X"00",
41641=>X"00",
41642=>X"00",
41643=>X"00",
41644=>X"00",
41645=>X"00",
41646=>X"00",
41647=>X"00",
41648=>X"00",
41649=>X"00",
41650=>X"00",
41651=>X"00",
41652=>X"00",
41653=>X"00",
41654=>X"00",
41655=>X"00",
41656=>X"00",
41657=>X"00",
41658=>X"00",
41659=>X"00",
41660=>X"00",
41661=>X"00",
41662=>X"00",
41663=>X"00",
41664=>X"00",
41665=>X"00",
41666=>X"00",
41667=>X"00",
41668=>X"00",
41669=>X"00",
41670=>X"00",
41671=>X"00",
41672=>X"00",
41673=>X"00",
41674=>X"00",
41675=>X"00",
41676=>X"00",
41677=>X"00",
41678=>X"00",
41679=>X"00",
41680=>X"00",
41681=>X"00",
41682=>X"00",
41683=>X"00",
41684=>X"00",
41685=>X"00",
41686=>X"00",
41687=>X"00",
41688=>X"00",
41689=>X"00",
41690=>X"00",
41691=>X"00",
41692=>X"00",
41693=>X"00",
41694=>X"00",
41695=>X"00",
41696=>X"00",
41697=>X"00",
41698=>X"00",
41699=>X"00",
41700=>X"00",
41701=>X"00",
41702=>X"00",
41703=>X"00",
41704=>X"00",
41705=>X"00",
41706=>X"00",
41707=>X"00",
41708=>X"00",
41709=>X"00",
41710=>X"00",
41711=>X"00",
41712=>X"00",
41713=>X"00",
41714=>X"00",
41715=>X"00",
41716=>X"00",
41717=>X"00",
41718=>X"00",
41719=>X"00",
41720=>X"00",
41721=>X"00",
41722=>X"00",
41723=>X"00",
41724=>X"00",
41725=>X"00",
41726=>X"00",
41727=>X"00",
41728=>X"00",
41729=>X"00",
41730=>X"00",
41731=>X"00",
41732=>X"00",
41733=>X"00",
41734=>X"00",
41735=>X"00",
41736=>X"00",
41737=>X"00",
41738=>X"00",
41739=>X"00",
41740=>X"00",
41741=>X"00",
41742=>X"00",
41743=>X"00",
41744=>X"00",
41745=>X"00",
41746=>X"00",
41747=>X"00",
41748=>X"00",
41749=>X"00",
41750=>X"00",
41751=>X"00",
41752=>X"00",
41753=>X"00",
41754=>X"00",
41755=>X"00",
41756=>X"00",
41757=>X"00",
41758=>X"00",
41759=>X"00",
41760=>X"00",
41761=>X"00",
41762=>X"00",
41763=>X"00",
41764=>X"00",
41765=>X"00",
41766=>X"00",
41767=>X"00",
41768=>X"00",
41769=>X"00",
41770=>X"00",
41771=>X"00",
41772=>X"00",
41773=>X"00",
41774=>X"00",
41775=>X"00",
41776=>X"00",
41777=>X"00",
41778=>X"00",
41779=>X"00",
41780=>X"00",
41781=>X"00",
41782=>X"00",
41783=>X"00",
41784=>X"00",
41785=>X"00",
41786=>X"00",
41787=>X"00",
41788=>X"00",
41789=>X"00",
41790=>X"00",
41791=>X"00",
41792=>X"00",
41793=>X"00",
41794=>X"00",
41795=>X"00",
41796=>X"00",
41797=>X"00",
41798=>X"00",
41799=>X"00",
41800=>X"00",
41801=>X"00",
41802=>X"00",
41803=>X"00",
41804=>X"00",
41805=>X"00",
41806=>X"00",
41807=>X"00",
41808=>X"00",
41809=>X"00",
41810=>X"00",
41811=>X"00",
41812=>X"00",
41813=>X"00",
41814=>X"00",
41815=>X"00",
41816=>X"00",
41817=>X"00",
41818=>X"00",
41819=>X"00",
41820=>X"00",
41821=>X"00",
41822=>X"00",
41823=>X"00",
41824=>X"00",
41825=>X"00",
41826=>X"00",
41827=>X"00",
41828=>X"00",
41829=>X"00",
41830=>X"00",
41831=>X"00",
41832=>X"00",
41833=>X"00",
41834=>X"00",
41835=>X"00",
41836=>X"00",
41837=>X"00",
41838=>X"00",
41839=>X"00",
41840=>X"00",
41841=>X"00",
41842=>X"00",
41843=>X"00",
41844=>X"00",
41845=>X"00",
41846=>X"00",
41847=>X"00",
41848=>X"00",
41849=>X"00",
41850=>X"00",
41851=>X"00",
41852=>X"00",
41853=>X"00",
41854=>X"00",
41855=>X"00",
41856=>X"00",
41857=>X"00",
41858=>X"00",
41859=>X"00",
41860=>X"00",
41861=>X"00",
41862=>X"00",
41863=>X"00",
41864=>X"00",
41865=>X"00",
41866=>X"00",
41867=>X"00",
41868=>X"00",
41869=>X"00",
41870=>X"00",
41871=>X"00",
41872=>X"00",
41873=>X"00",
41874=>X"00",
41875=>X"00",
41876=>X"00",
41877=>X"00",
41878=>X"00",
41879=>X"00",
41880=>X"00",
41881=>X"00",
41882=>X"00",
41883=>X"00",
41884=>X"00",
41885=>X"00",
41886=>X"00",
41887=>X"00",
41888=>X"00",
41889=>X"00",
41890=>X"00",
41891=>X"00",
41892=>X"00",
41893=>X"00",
41894=>X"00",
41895=>X"00",
41896=>X"00",
41897=>X"00",
41898=>X"00",
41899=>X"00",
41900=>X"00",
41901=>X"00",
41902=>X"00",
41903=>X"00",
41904=>X"00",
41905=>X"00",
41906=>X"00",
41907=>X"00",
41908=>X"00",
41909=>X"00",
41910=>X"00",
41911=>X"00",
41912=>X"00",
41913=>X"00",
41914=>X"00",
41915=>X"00",
41916=>X"00",
41917=>X"00",
41918=>X"00",
41919=>X"00",
41920=>X"00",
41921=>X"00",
41922=>X"00",
41923=>X"00",
41924=>X"00",
41925=>X"00",
41926=>X"00",
41927=>X"00",
41928=>X"00",
41929=>X"00",
41930=>X"00",
41931=>X"00",
41932=>X"00",
41933=>X"00",
41934=>X"00",
41935=>X"00",
41936=>X"00",
41937=>X"00",
41938=>X"00",
41939=>X"00",
41940=>X"00",
41941=>X"00",
41942=>X"00",
41943=>X"00",
41944=>X"00",
41945=>X"00",
41946=>X"00",
41947=>X"00",
41948=>X"00",
41949=>X"00",
41950=>X"00",
41951=>X"00",
41952=>X"00",
41953=>X"00",
41954=>X"00",
41955=>X"00",
41956=>X"00",
41957=>X"00",
41958=>X"00",
41959=>X"00",
41960=>X"00",
41961=>X"00",
41962=>X"00",
41963=>X"00",
41964=>X"00",
41965=>X"00",
41966=>X"00",
41967=>X"00",
41968=>X"00",
41969=>X"00",
41970=>X"00",
41971=>X"00",
41972=>X"00",
41973=>X"00",
41974=>X"00",
41975=>X"00",
41976=>X"00",
41977=>X"00",
41978=>X"00",
41979=>X"00",
41980=>X"00",
41981=>X"00",
41982=>X"00",
41983=>X"00",
41984=>X"00",
41985=>X"00",
41986=>X"00",
41987=>X"00",
41988=>X"00",
41989=>X"00",
41990=>X"00",
41991=>X"00",
41992=>X"00",
41993=>X"00",
41994=>X"00",
41995=>X"00",
41996=>X"00",
41997=>X"00",
41998=>X"00",
41999=>X"00",
42000=>X"00",
42001=>X"00",
42002=>X"00",
42003=>X"00",
42004=>X"00",
42005=>X"00",
42006=>X"00",
42007=>X"00",
42008=>X"00",
42009=>X"00",
42010=>X"00",
42011=>X"00",
42012=>X"00",
42013=>X"00",
42014=>X"00",
42015=>X"00",
42016=>X"00",
42017=>X"00",
42018=>X"00",
42019=>X"00",
42020=>X"00",
42021=>X"00",
42022=>X"00",
42023=>X"00",
42024=>X"00",
42025=>X"00",
42026=>X"00",
42027=>X"00",
42028=>X"00",
42029=>X"00",
42030=>X"00",
42031=>X"00",
42032=>X"00",
42033=>X"00",
42034=>X"00",
42035=>X"00",
42036=>X"00",
42037=>X"00",
42038=>X"00",
42039=>X"00",
42040=>X"00",
42041=>X"00",
42042=>X"00",
42043=>X"00",
42044=>X"00",
42045=>X"00",
42046=>X"00",
42047=>X"00",
42048=>X"00",
42049=>X"00",
42050=>X"00",
42051=>X"00",
42052=>X"00",
42053=>X"00",
42054=>X"00",
42055=>X"00",
42056=>X"00",
42057=>X"00",
42058=>X"00",
42059=>X"00",
42060=>X"00",
42061=>X"00",
42062=>X"00",
42063=>X"00",
42064=>X"00",
42065=>X"00",
42066=>X"00",
42067=>X"00",
42068=>X"00",
42069=>X"00",
42070=>X"00",
42071=>X"00",
42072=>X"00",
42073=>X"00",
42074=>X"00",
42075=>X"00",
42076=>X"00",
42077=>X"00",
42078=>X"00",
42079=>X"00",
42080=>X"00",
42081=>X"00",
42082=>X"00",
42083=>X"00",
42084=>X"00",
42085=>X"00",
42086=>X"00",
42087=>X"00",
42088=>X"00",
42089=>X"00",
42090=>X"00",
42091=>X"00",
42092=>X"00",
42093=>X"00",
42094=>X"00",
42095=>X"00",
42096=>X"00",
42097=>X"00",
42098=>X"00",
42099=>X"00",
42100=>X"00",
42101=>X"00",
42102=>X"00",
42103=>X"00",
42104=>X"00",
42105=>X"00",
42106=>X"00",
42107=>X"00",
42108=>X"00",
42109=>X"00",
42110=>X"00",
42111=>X"00",
42112=>X"00",
42113=>X"00",
42114=>X"00",
42115=>X"00",
42116=>X"00",
42117=>X"00",
42118=>X"00",
42119=>X"00",
42120=>X"00",
42121=>X"00",
42122=>X"00",
42123=>X"00",
42124=>X"00",
42125=>X"00",
42126=>X"00",
42127=>X"00",
42128=>X"00",
42129=>X"00",
42130=>X"00",
42131=>X"00",
42132=>X"00",
42133=>X"00",
42134=>X"00",
42135=>X"00",
42136=>X"00",
42137=>X"00",
42138=>X"00",
42139=>X"00",
42140=>X"00",
42141=>X"00",
42142=>X"00",
42143=>X"00",
42144=>X"00",
42145=>X"00",
42146=>X"00",
42147=>X"00",
42148=>X"00",
42149=>X"00",
42150=>X"00",
42151=>X"00",
42152=>X"00",
42153=>X"00",
42154=>X"00",
42155=>X"00",
42156=>X"00",
42157=>X"00",
42158=>X"00",
42159=>X"00",
42160=>X"00",
42161=>X"00",
42162=>X"00",
42163=>X"00",
42164=>X"00",
42165=>X"00",
42166=>X"00",
42167=>X"00",
42168=>X"00",
42169=>X"00",
42170=>X"00",
42171=>X"00",
42172=>X"00",
42173=>X"00",
42174=>X"00",
42175=>X"00",
42176=>X"00",
42177=>X"00",
42178=>X"00",
42179=>X"00",
42180=>X"00",
42181=>X"00",
42182=>X"00",
42183=>X"00",
42184=>X"00",
42185=>X"00",
42186=>X"00",
42187=>X"00",
42188=>X"00",
42189=>X"00",
42190=>X"00",
42191=>X"00",
42192=>X"00",
42193=>X"00",
42194=>X"00",
42195=>X"00",
42196=>X"00",
42197=>X"00",
42198=>X"00",
42199=>X"00",
42200=>X"00",
42201=>X"00",
42202=>X"00",
42203=>X"00",
42204=>X"00",
42205=>X"00",
42206=>X"00",
42207=>X"00",
42208=>X"00",
42209=>X"00",
42210=>X"00",
42211=>X"00",
42212=>X"00",
42213=>X"00",
42214=>X"00",
42215=>X"00",
42216=>X"00",
42217=>X"00",
42218=>X"00",
42219=>X"00",
42220=>X"00",
42221=>X"00",
42222=>X"00",
42223=>X"00",
42224=>X"00",
42225=>X"00",
42226=>X"00",
42227=>X"00",
42228=>X"00",
42229=>X"00",
42230=>X"00",
42231=>X"00",
42232=>X"00",
42233=>X"00",
42234=>X"00",
42235=>X"00",
42236=>X"00",
42237=>X"00",
42238=>X"00",
42239=>X"00",
42240=>X"00",
42241=>X"00",
42242=>X"00",
42243=>X"00",
42244=>X"00",
42245=>X"00",
42246=>X"00",
42247=>X"00",
42248=>X"00",
42249=>X"00",
42250=>X"00",
42251=>X"00",
42252=>X"00",
42253=>X"00",
42254=>X"00",
42255=>X"00",
42256=>X"00",
42257=>X"00",
42258=>X"00",
42259=>X"00",
42260=>X"00",
42261=>X"00",
42262=>X"00",
42263=>X"00",
42264=>X"00",
42265=>X"00",
42266=>X"00",
42267=>X"00",
42268=>X"00",
42269=>X"00",
42270=>X"00",
42271=>X"00",
42272=>X"00",
42273=>X"00",
42274=>X"00",
42275=>X"00",
42276=>X"00",
42277=>X"00",
42278=>X"00",
42279=>X"00",
42280=>X"00",
42281=>X"00",
42282=>X"00",
42283=>X"00",
42284=>X"00",
42285=>X"00",
42286=>X"00",
42287=>X"00",
42288=>X"00",
42289=>X"00",
42290=>X"00",
42291=>X"00",
42292=>X"00",
42293=>X"00",
42294=>X"00",
42295=>X"00",
42296=>X"00",
42297=>X"00",
42298=>X"00",
42299=>X"00",
42300=>X"00",
42301=>X"00",
42302=>X"00",
42303=>X"00",
42304=>X"00",
42305=>X"00",
42306=>X"00",
42307=>X"00",
42308=>X"00",
42309=>X"00",
42310=>X"00",
42311=>X"00",
42312=>X"00",
42313=>X"00",
42314=>X"00",
42315=>X"00",
42316=>X"00",
42317=>X"00",
42318=>X"00",
42319=>X"00",
42320=>X"00",
42321=>X"00",
42322=>X"00",
42323=>X"00",
42324=>X"00",
42325=>X"00",
42326=>X"00",
42327=>X"00",
42328=>X"00",
42329=>X"00",
42330=>X"00",
42331=>X"00",
42332=>X"00",
42333=>X"00",
42334=>X"00",
42335=>X"00",
42336=>X"00",
42337=>X"00",
42338=>X"00",
42339=>X"00",
42340=>X"00",
42341=>X"00",
42342=>X"00",
42343=>X"00",
42344=>X"00",
42345=>X"00",
42346=>X"00",
42347=>X"00",
42348=>X"00",
42349=>X"00",
42350=>X"00",
42351=>X"00",
42352=>X"00",
42353=>X"00",
42354=>X"00",
42355=>X"00",
42356=>X"00",
42357=>X"00",
42358=>X"00",
42359=>X"00",
42360=>X"00",
42361=>X"00",
42362=>X"00",
42363=>X"00",
42364=>X"00",
42365=>X"00",
42366=>X"00",
42367=>X"00",
42368=>X"00",
42369=>X"00",
42370=>X"00",
42371=>X"00",
42372=>X"00",
42373=>X"00",
42374=>X"00",
42375=>X"00",
42376=>X"00",
42377=>X"00",
42378=>X"00",
42379=>X"00",
42380=>X"00",
42381=>X"00",
42382=>X"00",
42383=>X"00",
42384=>X"00",
42385=>X"00",
42386=>X"00",
42387=>X"00",
42388=>X"00",
42389=>X"00",
42390=>X"00",
42391=>X"00",
42392=>X"00",
42393=>X"00",
42394=>X"00",
42395=>X"00",
42396=>X"00",
42397=>X"00",
42398=>X"00",
42399=>X"00",
42400=>X"00",
42401=>X"00",
42402=>X"00",
42403=>X"00",
42404=>X"00",
42405=>X"00",
42406=>X"00",
42407=>X"00",
42408=>X"00",
42409=>X"00",
42410=>X"00",
42411=>X"00",
42412=>X"00",
42413=>X"00",
42414=>X"00",
42415=>X"00",
42416=>X"00",
42417=>X"00",
42418=>X"00",
42419=>X"00",
42420=>X"00",
42421=>X"00",
42422=>X"00",
42423=>X"00",
42424=>X"00",
42425=>X"00",
42426=>X"00",
42427=>X"00",
42428=>X"00",
42429=>X"00",
42430=>X"00",
42431=>X"00",
42432=>X"00",
42433=>X"00",
42434=>X"00",
42435=>X"00",
42436=>X"00",
42437=>X"00",
42438=>X"00",
42439=>X"00",
42440=>X"00",
42441=>X"00",
42442=>X"00",
42443=>X"00",
42444=>X"00",
42445=>X"00",
42446=>X"00",
42447=>X"00",
42448=>X"00",
42449=>X"00",
42450=>X"00",
42451=>X"00",
42452=>X"00",
42453=>X"00",
42454=>X"00",
42455=>X"00",
42456=>X"00",
42457=>X"00",
42458=>X"00",
42459=>X"00",
42460=>X"00",
42461=>X"00",
42462=>X"00",
42463=>X"00",
42464=>X"00",
42465=>X"00",
42466=>X"00",
42467=>X"00",
42468=>X"00",
42469=>X"00",
42470=>X"00",
42471=>X"00",
42472=>X"00",
42473=>X"00",
42474=>X"00",
42475=>X"00",
42476=>X"00",
42477=>X"00",
42478=>X"00",
42479=>X"00",
42480=>X"00",
42481=>X"00",
42482=>X"00",
42483=>X"00",
42484=>X"00",
42485=>X"00",
42486=>X"00",
42487=>X"00",
42488=>X"00",
42489=>X"00",
42490=>X"00",
42491=>X"00",
42492=>X"00",
42493=>X"00",
42494=>X"00",
42495=>X"00",
42496=>X"00",
42497=>X"00",
42498=>X"00",
42499=>X"00",
42500=>X"00",
42501=>X"00",
42502=>X"00",
42503=>X"00",
42504=>X"00",
42505=>X"00",
42506=>X"00",
42507=>X"00",
42508=>X"00",
42509=>X"00",
42510=>X"00",
42511=>X"00",
42512=>X"00",
42513=>X"00",
42514=>X"00",
42515=>X"00",
42516=>X"00",
42517=>X"00",
42518=>X"00",
42519=>X"00",
42520=>X"00",
42521=>X"00",
42522=>X"00",
42523=>X"00",
42524=>X"00",
42525=>X"00",
42526=>X"00",
42527=>X"00",
42528=>X"00",
42529=>X"00",
42530=>X"00",
42531=>X"00",
42532=>X"00",
42533=>X"00",
42534=>X"00",
42535=>X"00",
42536=>X"00",
42537=>X"00",
42538=>X"00",
42539=>X"00",
42540=>X"00",
42541=>X"00",
42542=>X"00",
42543=>X"00",
42544=>X"00",
42545=>X"00",
42546=>X"00",
42547=>X"00",
42548=>X"00",
42549=>X"00",
42550=>X"00",
42551=>X"00",
42552=>X"00",
42553=>X"00",
42554=>X"00",
42555=>X"00",
42556=>X"00",
42557=>X"00",
42558=>X"00",
42559=>X"00",
42560=>X"00",
42561=>X"00",
42562=>X"00",
42563=>X"00",
42564=>X"00",
42565=>X"00",
42566=>X"00",
42567=>X"00",
42568=>X"00",
42569=>X"00",
42570=>X"00",
42571=>X"00",
42572=>X"00",
42573=>X"00",
42574=>X"00",
42575=>X"00",
42576=>X"00",
42577=>X"00",
42578=>X"00",
42579=>X"00",
42580=>X"00",
42581=>X"00",
42582=>X"00",
42583=>X"00",
42584=>X"00",
42585=>X"00",
42586=>X"00",
42587=>X"00",
42588=>X"00",
42589=>X"00",
42590=>X"00",
42591=>X"00",
42592=>X"00",
42593=>X"00",
42594=>X"00",
42595=>X"00",
42596=>X"00",
42597=>X"00",
42598=>X"00",
42599=>X"00",
42600=>X"00",
42601=>X"00",
42602=>X"00",
42603=>X"00",
42604=>X"00",
42605=>X"00",
42606=>X"00",
42607=>X"00",
42608=>X"00",
42609=>X"00",
42610=>X"00",
42611=>X"00",
42612=>X"00",
42613=>X"00",
42614=>X"00",
42615=>X"00",
42616=>X"00",
42617=>X"00",
42618=>X"00",
42619=>X"00",
42620=>X"00",
42621=>X"00",
42622=>X"00",
42623=>X"00",
42624=>X"00",
42625=>X"00",
42626=>X"00",
42627=>X"00",
42628=>X"00",
42629=>X"00",
42630=>X"00",
42631=>X"00",
42632=>X"00",
42633=>X"00",
42634=>X"00",
42635=>X"00",
42636=>X"00",
42637=>X"00",
42638=>X"00",
42639=>X"00",
42640=>X"00",
42641=>X"00",
42642=>X"00",
42643=>X"00",
42644=>X"00",
42645=>X"00",
42646=>X"00",
42647=>X"00",
42648=>X"00",
42649=>X"00",
42650=>X"00",
42651=>X"00",
42652=>X"00",
42653=>X"00",
42654=>X"00",
42655=>X"00",
42656=>X"00",
42657=>X"00",
42658=>X"00",
42659=>X"00",
42660=>X"00",
42661=>X"00",
42662=>X"00",
42663=>X"00",
42664=>X"00",
42665=>X"00",
42666=>X"00",
42667=>X"00",
42668=>X"00",
42669=>X"00",
42670=>X"00",
42671=>X"00",
42672=>X"00",
42673=>X"00",
42674=>X"00",
42675=>X"00",
42676=>X"00",
42677=>X"00",
42678=>X"00",
42679=>X"00",
42680=>X"00",
42681=>X"00",
42682=>X"00",
42683=>X"00",
42684=>X"00",
42685=>X"00",
42686=>X"00",
42687=>X"00",
42688=>X"00",
42689=>X"00",
42690=>X"00",
42691=>X"00",
42692=>X"00",
42693=>X"00",
42694=>X"00",
42695=>X"00",
42696=>X"00",
42697=>X"00",
42698=>X"00",
42699=>X"00",
42700=>X"00",
42701=>X"00",
42702=>X"00",
42703=>X"00",
42704=>X"00",
42705=>X"00",
42706=>X"00",
42707=>X"00",
42708=>X"00",
42709=>X"00",
42710=>X"00",
42711=>X"00",
42712=>X"00",
42713=>X"00",
42714=>X"00",
42715=>X"00",
42716=>X"00",
42717=>X"00",
42718=>X"00",
42719=>X"00",
42720=>X"00",
42721=>X"00",
42722=>X"00",
42723=>X"00",
42724=>X"00",
42725=>X"00",
42726=>X"00",
42727=>X"00",
42728=>X"00",
42729=>X"00",
42730=>X"00",
42731=>X"00",
42732=>X"00",
42733=>X"00",
42734=>X"00",
42735=>X"00",
42736=>X"00",
42737=>X"00",
42738=>X"00",
42739=>X"00",
42740=>X"00",
42741=>X"00",
42742=>X"00",
42743=>X"00",
42744=>X"00",
42745=>X"00",
42746=>X"00",
42747=>X"00",
42748=>X"00",
42749=>X"00",
42750=>X"00",
42751=>X"00",
42752=>X"00",
42753=>X"00",
42754=>X"00",
42755=>X"00",
42756=>X"00",
42757=>X"00",
42758=>X"00",
42759=>X"00",
42760=>X"00",
42761=>X"00",
42762=>X"00",
42763=>X"00",
42764=>X"00",
42765=>X"00",
42766=>X"00",
42767=>X"00",
42768=>X"00",
42769=>X"00",
42770=>X"00",
42771=>X"00",
42772=>X"00",
42773=>X"00",
42774=>X"00",
42775=>X"00",
42776=>X"00",
42777=>X"00",
42778=>X"00",
42779=>X"00",
42780=>X"00",
42781=>X"00",
42782=>X"00",
42783=>X"00",
42784=>X"00",
42785=>X"00",
42786=>X"00",
42787=>X"00",
42788=>X"00",
42789=>X"00",
42790=>X"00",
42791=>X"00",
42792=>X"00",
42793=>X"00",
42794=>X"00",
42795=>X"00",
42796=>X"00",
42797=>X"00",
42798=>X"00",
42799=>X"00",
42800=>X"00",
42801=>X"00",
42802=>X"00",
42803=>X"00",
42804=>X"00",
42805=>X"00",
42806=>X"00",
42807=>X"00",
42808=>X"00",
42809=>X"00",
42810=>X"00",
42811=>X"00",
42812=>X"00",
42813=>X"00",
42814=>X"00",
42815=>X"00",
42816=>X"00",
42817=>X"00",
42818=>X"00",
42819=>X"00",
42820=>X"00",
42821=>X"00",
42822=>X"00",
42823=>X"00",
42824=>X"00",
42825=>X"00",
42826=>X"00",
42827=>X"00",
42828=>X"00",
42829=>X"00",
42830=>X"00",
42831=>X"00",
42832=>X"00",
42833=>X"00",
42834=>X"00",
42835=>X"00",
42836=>X"00",
42837=>X"00",
42838=>X"00",
42839=>X"00",
42840=>X"00",
42841=>X"00",
42842=>X"00",
42843=>X"00",
42844=>X"00",
42845=>X"00",
42846=>X"00",
42847=>X"00",
42848=>X"00",
42849=>X"00",
42850=>X"00",
42851=>X"00",
42852=>X"00",
42853=>X"00",
42854=>X"00",
42855=>X"00",
42856=>X"00",
42857=>X"00",
42858=>X"00",
42859=>X"00",
42860=>X"00",
42861=>X"00",
42862=>X"00",
42863=>X"00",
42864=>X"00",
42865=>X"00",
42866=>X"00",
42867=>X"00",
42868=>X"00",
42869=>X"00",
42870=>X"00",
42871=>X"00",
42872=>X"00",
42873=>X"00",
42874=>X"00",
42875=>X"00",
42876=>X"00",
42877=>X"00",
42878=>X"00",
42879=>X"00",
42880=>X"00",
42881=>X"00",
42882=>X"00",
42883=>X"00",
42884=>X"00",
42885=>X"00",
42886=>X"00",
42887=>X"00",
42888=>X"00",
42889=>X"00",
42890=>X"00",
42891=>X"00",
42892=>X"00",
42893=>X"00",
42894=>X"00",
42895=>X"00",
42896=>X"00",
42897=>X"00",
42898=>X"00",
42899=>X"00",
42900=>X"00",
42901=>X"00",
42902=>X"00",
42903=>X"00",
42904=>X"00",
42905=>X"00",
42906=>X"00",
42907=>X"00",
42908=>X"00",
42909=>X"00",
42910=>X"00",
42911=>X"00",
42912=>X"00",
42913=>X"00",
42914=>X"00",
42915=>X"00",
42916=>X"00",
42917=>X"00",
42918=>X"00",
42919=>X"00",
42920=>X"00",
42921=>X"00",
42922=>X"00",
42923=>X"00",
42924=>X"00",
42925=>X"00",
42926=>X"00",
42927=>X"00",
42928=>X"00",
42929=>X"00",
42930=>X"00",
42931=>X"00",
42932=>X"00",
42933=>X"00",
42934=>X"00",
42935=>X"00",
42936=>X"00",
42937=>X"00",
42938=>X"00",
42939=>X"00",
42940=>X"00",
42941=>X"00",
42942=>X"00",
42943=>X"00",
42944=>X"00",
42945=>X"00",
42946=>X"00",
42947=>X"00",
42948=>X"00",
42949=>X"00",
42950=>X"00",
42951=>X"00",
42952=>X"00",
42953=>X"00",
42954=>X"00",
42955=>X"00",
42956=>X"00",
42957=>X"00",
42958=>X"00",
42959=>X"00",
42960=>X"00",
42961=>X"00",
42962=>X"00",
42963=>X"00",
42964=>X"00",
42965=>X"00",
42966=>X"00",
42967=>X"00",
42968=>X"00",
42969=>X"00",
42970=>X"00",
42971=>X"00",
42972=>X"00",
42973=>X"00",
42974=>X"00",
42975=>X"00",
42976=>X"00",
42977=>X"00",
42978=>X"00",
42979=>X"00",
42980=>X"00",
42981=>X"00",
42982=>X"00",
42983=>X"00",
42984=>X"00",
42985=>X"00",
42986=>X"00",
42987=>X"00",
42988=>X"00",
42989=>X"00",
42990=>X"00",
42991=>X"00",
42992=>X"00",
42993=>X"00",
42994=>X"00",
42995=>X"00",
42996=>X"00",
42997=>X"00",
42998=>X"00",
42999=>X"00",
43000=>X"00",
43001=>X"00",
43002=>X"00",
43003=>X"00",
43004=>X"00",
43005=>X"00",
43006=>X"00",
43007=>X"00",
43008=>X"00",
43009=>X"00",
43010=>X"00",
43011=>X"00",
43012=>X"00",
43013=>X"00",
43014=>X"00",
43015=>X"00",
43016=>X"00",
43017=>X"00",
43018=>X"00",
43019=>X"00",
43020=>X"00",
43021=>X"00",
43022=>X"00",
43023=>X"00",
43024=>X"00",
43025=>X"00",
43026=>X"00",
43027=>X"00",
43028=>X"00",
43029=>X"00",
43030=>X"00",
43031=>X"00",
43032=>X"00",
43033=>X"00",
43034=>X"00",
43035=>X"00",
43036=>X"00",
43037=>X"00",
43038=>X"00",
43039=>X"00",
43040=>X"00",
43041=>X"00",
43042=>X"00",
43043=>X"00",
43044=>X"00",
43045=>X"00",
43046=>X"00",
43047=>X"00",
43048=>X"00",
43049=>X"00",
43050=>X"00",
43051=>X"00",
43052=>X"00",
43053=>X"00",
43054=>X"00",
43055=>X"00",
43056=>X"00",
43057=>X"00",
43058=>X"00",
43059=>X"00",
43060=>X"00",
43061=>X"00",
43062=>X"00",
43063=>X"00",
43064=>X"00",
43065=>X"00",
43066=>X"00",
43067=>X"00",
43068=>X"00",
43069=>X"00",
43070=>X"00",
43071=>X"00",
43072=>X"00",
43073=>X"00",
43074=>X"00",
43075=>X"00",
43076=>X"00",
43077=>X"00",
43078=>X"00",
43079=>X"00",
43080=>X"00",
43081=>X"00",
43082=>X"00",
43083=>X"00",
43084=>X"00",
43085=>X"00",
43086=>X"00",
43087=>X"00",
43088=>X"00",
43089=>X"00",
43090=>X"00",
43091=>X"00",
43092=>X"00",
43093=>X"00",
43094=>X"00",
43095=>X"00",
43096=>X"00",
43097=>X"00",
43098=>X"00",
43099=>X"00",
43100=>X"00",
43101=>X"00",
43102=>X"00",
43103=>X"00",
43104=>X"00",
43105=>X"00",
43106=>X"00",
43107=>X"00",
43108=>X"00",
43109=>X"00",
43110=>X"00",
43111=>X"00",
43112=>X"00",
43113=>X"00",
43114=>X"00",
43115=>X"00",
43116=>X"00",
43117=>X"00",
43118=>X"00",
43119=>X"00",
43120=>X"00",
43121=>X"00",
43122=>X"00",
43123=>X"00",
43124=>X"00",
43125=>X"00",
43126=>X"00",
43127=>X"00",
43128=>X"00",
43129=>X"00",
43130=>X"00",
43131=>X"00",
43132=>X"00",
43133=>X"00",
43134=>X"00",
43135=>X"00",
43136=>X"00",
43137=>X"00",
43138=>X"00",
43139=>X"00",
43140=>X"00",
43141=>X"00",
43142=>X"00",
43143=>X"00",
43144=>X"00",
43145=>X"00",
43146=>X"00",
43147=>X"00",
43148=>X"00",
43149=>X"00",
43150=>X"00",
43151=>X"00",
43152=>X"00",
43153=>X"00",
43154=>X"00",
43155=>X"00",
43156=>X"00",
43157=>X"00",
43158=>X"00",
43159=>X"00",
43160=>X"00",
43161=>X"00",
43162=>X"00",
43163=>X"00",
43164=>X"00",
43165=>X"00",
43166=>X"00",
43167=>X"00",
43168=>X"00",
43169=>X"00",
43170=>X"00",
43171=>X"00",
43172=>X"00",
43173=>X"00",
43174=>X"00",
43175=>X"00",
43176=>X"00",
43177=>X"00",
43178=>X"00",
43179=>X"00",
43180=>X"00",
43181=>X"00",
43182=>X"00",
43183=>X"00",
43184=>X"00",
43185=>X"00",
43186=>X"00",
43187=>X"00",
43188=>X"00",
43189=>X"00",
43190=>X"00",
43191=>X"00",
43192=>X"00",
43193=>X"00",
43194=>X"00",
43195=>X"00",
43196=>X"00",
43197=>X"00",
43198=>X"00",
43199=>X"00",
43200=>X"00",
43201=>X"00",
43202=>X"00",
43203=>X"00",
43204=>X"00",
43205=>X"00",
43206=>X"00",
43207=>X"00",
43208=>X"00",
43209=>X"00",
43210=>X"00",
43211=>X"00",
43212=>X"00",
43213=>X"00",
43214=>X"00",
43215=>X"00",
43216=>X"00",
43217=>X"00",
43218=>X"00",
43219=>X"00",
43220=>X"00",
43221=>X"00",
43222=>X"00",
43223=>X"00",
43224=>X"00",
43225=>X"00",
43226=>X"00",
43227=>X"00",
43228=>X"00",
43229=>X"00",
43230=>X"00",
43231=>X"00",
43232=>X"00",
43233=>X"00",
43234=>X"00",
43235=>X"00",
43236=>X"00",
43237=>X"00",
43238=>X"00",
43239=>X"00",
43240=>X"00",
43241=>X"00",
43242=>X"00",
43243=>X"00",
43244=>X"00",
43245=>X"00",
43246=>X"00",
43247=>X"00",
43248=>X"00",
43249=>X"00",
43250=>X"00",
43251=>X"00",
43252=>X"00",
43253=>X"00",
43254=>X"00",
43255=>X"00",
43256=>X"00",
43257=>X"00",
43258=>X"00",
43259=>X"00",
43260=>X"00",
43261=>X"00",
43262=>X"00",
43263=>X"00",
43264=>X"00",
43265=>X"00",
43266=>X"00",
43267=>X"00",
43268=>X"00",
43269=>X"00",
43270=>X"00",
43271=>X"00",
43272=>X"00",
43273=>X"00",
43274=>X"00",
43275=>X"00",
43276=>X"00",
43277=>X"00",
43278=>X"00",
43279=>X"00",
43280=>X"00",
43281=>X"00",
43282=>X"00",
43283=>X"00",
43284=>X"00",
43285=>X"00",
43286=>X"00",
43287=>X"00",
43288=>X"00",
43289=>X"00",
43290=>X"00",
43291=>X"00",
43292=>X"00",
43293=>X"00",
43294=>X"00",
43295=>X"00",
43296=>X"00",
43297=>X"00",
43298=>X"00",
43299=>X"00",
43300=>X"00",
43301=>X"00",
43302=>X"00",
43303=>X"00",
43304=>X"00",
43305=>X"00",
43306=>X"00",
43307=>X"00",
43308=>X"00",
43309=>X"00",
43310=>X"00",
43311=>X"00",
43312=>X"00",
43313=>X"00",
43314=>X"00",
43315=>X"00",
43316=>X"00",
43317=>X"00",
43318=>X"00",
43319=>X"00",
43320=>X"00",
43321=>X"00",
43322=>X"00",
43323=>X"00",
43324=>X"00",
43325=>X"00",
43326=>X"00",
43327=>X"00",
43328=>X"00",
43329=>X"00",
43330=>X"00",
43331=>X"00",
43332=>X"00",
43333=>X"00",
43334=>X"00",
43335=>X"00",
43336=>X"00",
43337=>X"00",
43338=>X"00",
43339=>X"00",
43340=>X"00",
43341=>X"00",
43342=>X"00",
43343=>X"00",
43344=>X"00",
43345=>X"00",
43346=>X"00",
43347=>X"00",
43348=>X"00",
43349=>X"00",
43350=>X"00",
43351=>X"00",
43352=>X"00",
43353=>X"00",
43354=>X"00",
43355=>X"00",
43356=>X"00",
43357=>X"00",
43358=>X"00",
43359=>X"00",
43360=>X"00",
43361=>X"00",
43362=>X"00",
43363=>X"00",
43364=>X"00",
43365=>X"00",
43366=>X"00",
43367=>X"00",
43368=>X"00",
43369=>X"00",
43370=>X"00",
43371=>X"00",
43372=>X"00",
43373=>X"00",
43374=>X"00",
43375=>X"00",
43376=>X"00",
43377=>X"00",
43378=>X"00",
43379=>X"00",
43380=>X"00",
43381=>X"00",
43382=>X"00",
43383=>X"00",
43384=>X"00",
43385=>X"00",
43386=>X"00",
43387=>X"00",
43388=>X"00",
43389=>X"00",
43390=>X"00",
43391=>X"00",
43392=>X"00",
43393=>X"00",
43394=>X"00",
43395=>X"00",
43396=>X"00",
43397=>X"00",
43398=>X"00",
43399=>X"00",
43400=>X"00",
43401=>X"00",
43402=>X"00",
43403=>X"00",
43404=>X"00",
43405=>X"00",
43406=>X"00",
43407=>X"00",
43408=>X"00",
43409=>X"00",
43410=>X"00",
43411=>X"00",
43412=>X"00",
43413=>X"00",
43414=>X"00",
43415=>X"00",
43416=>X"00",
43417=>X"00",
43418=>X"00",
43419=>X"00",
43420=>X"00",
43421=>X"00",
43422=>X"00",
43423=>X"00",
43424=>X"00",
43425=>X"00",
43426=>X"00",
43427=>X"00",
43428=>X"00",
43429=>X"00",
43430=>X"00",
43431=>X"00",
43432=>X"00",
43433=>X"00",
43434=>X"00",
43435=>X"00",
43436=>X"00",
43437=>X"00",
43438=>X"00",
43439=>X"00",
43440=>X"00",
43441=>X"00",
43442=>X"00",
43443=>X"00",
43444=>X"00",
43445=>X"00",
43446=>X"00",
43447=>X"00",
43448=>X"00",
43449=>X"00",
43450=>X"00",
43451=>X"00",
43452=>X"00",
43453=>X"00",
43454=>X"00",
43455=>X"00",
43456=>X"00",
43457=>X"00",
43458=>X"00",
43459=>X"00",
43460=>X"00",
43461=>X"00",
43462=>X"00",
43463=>X"00",
43464=>X"00",
43465=>X"00",
43466=>X"00",
43467=>X"00",
43468=>X"00",
43469=>X"00",
43470=>X"00",
43471=>X"00",
43472=>X"00",
43473=>X"00",
43474=>X"00",
43475=>X"00",
43476=>X"00",
43477=>X"00",
43478=>X"00",
43479=>X"00",
43480=>X"00",
43481=>X"00",
43482=>X"00",
43483=>X"00",
43484=>X"00",
43485=>X"00",
43486=>X"00",
43487=>X"00",
43488=>X"00",
43489=>X"00",
43490=>X"00",
43491=>X"00",
43492=>X"00",
43493=>X"00",
43494=>X"00",
43495=>X"00",
43496=>X"00",
43497=>X"00",
43498=>X"00",
43499=>X"00",
43500=>X"00",
43501=>X"00",
43502=>X"00",
43503=>X"00",
43504=>X"00",
43505=>X"00",
43506=>X"00",
43507=>X"00",
43508=>X"00",
43509=>X"00",
43510=>X"00",
43511=>X"00",
43512=>X"00",
43513=>X"00",
43514=>X"00",
43515=>X"00",
43516=>X"00",
43517=>X"00",
43518=>X"00",
43519=>X"00",
43520=>X"00",
43521=>X"00",
43522=>X"00",
43523=>X"00",
43524=>X"00",
43525=>X"00",
43526=>X"00",
43527=>X"00",
43528=>X"00",
43529=>X"00",
43530=>X"00",
43531=>X"00",
43532=>X"00",
43533=>X"00",
43534=>X"00",
43535=>X"00",
43536=>X"00",
43537=>X"00",
43538=>X"00",
43539=>X"00",
43540=>X"00",
43541=>X"00",
43542=>X"00",
43543=>X"00",
43544=>X"00",
43545=>X"00",
43546=>X"00",
43547=>X"00",
43548=>X"00",
43549=>X"00",
43550=>X"00",
43551=>X"00",
43552=>X"00",
43553=>X"00",
43554=>X"00",
43555=>X"00",
43556=>X"00",
43557=>X"00",
43558=>X"00",
43559=>X"00",
43560=>X"00",
43561=>X"00",
43562=>X"00",
43563=>X"00",
43564=>X"00",
43565=>X"00",
43566=>X"00",
43567=>X"00",
43568=>X"00",
43569=>X"00",
43570=>X"00",
43571=>X"00",
43572=>X"00",
43573=>X"00",
43574=>X"00",
43575=>X"00",
43576=>X"00",
43577=>X"00",
43578=>X"00",
43579=>X"00",
43580=>X"00",
43581=>X"00",
43582=>X"00",
43583=>X"00",
43584=>X"00",
43585=>X"00",
43586=>X"00",
43587=>X"00",
43588=>X"00",
43589=>X"00",
43590=>X"00",
43591=>X"00",
43592=>X"00",
43593=>X"00",
43594=>X"00",
43595=>X"00",
43596=>X"00",
43597=>X"00",
43598=>X"00",
43599=>X"00",
43600=>X"00",
43601=>X"00",
43602=>X"00",
43603=>X"00",
43604=>X"00",
43605=>X"00",
43606=>X"00",
43607=>X"00",
43608=>X"00",
43609=>X"00",
43610=>X"00",
43611=>X"00",
43612=>X"00",
43613=>X"00",
43614=>X"00",
43615=>X"00",
43616=>X"00",
43617=>X"00",
43618=>X"00",
43619=>X"00",
43620=>X"00",
43621=>X"00",
43622=>X"00",
43623=>X"00",
43624=>X"00",
43625=>X"00",
43626=>X"00",
43627=>X"00",
43628=>X"00",
43629=>X"00",
43630=>X"00",
43631=>X"00",
43632=>X"00",
43633=>X"00",
43634=>X"00",
43635=>X"00",
43636=>X"00",
43637=>X"00",
43638=>X"00",
43639=>X"00",
43640=>X"00",
43641=>X"00",
43642=>X"00",
43643=>X"00",
43644=>X"00",
43645=>X"00",
43646=>X"00",
43647=>X"00",
43648=>X"00",
43649=>X"00",
43650=>X"00",
43651=>X"00",
43652=>X"00",
43653=>X"00",
43654=>X"00",
43655=>X"00",
43656=>X"00",
43657=>X"00",
43658=>X"00",
43659=>X"00",
43660=>X"00",
43661=>X"00",
43662=>X"00",
43663=>X"00",
43664=>X"00",
43665=>X"00",
43666=>X"00",
43667=>X"00",
43668=>X"00",
43669=>X"00",
43670=>X"00",
43671=>X"00",
43672=>X"00",
43673=>X"00",
43674=>X"00",
43675=>X"00",
43676=>X"00",
43677=>X"00",
43678=>X"00",
43679=>X"00",
43680=>X"00",
43681=>X"00",
43682=>X"00",
43683=>X"00",
43684=>X"00",
43685=>X"00",
43686=>X"00",
43687=>X"00",
43688=>X"00",
43689=>X"00",
43690=>X"00",
43691=>X"00",
43692=>X"00",
43693=>X"00",
43694=>X"00",
43695=>X"00",
43696=>X"00",
43697=>X"00",
43698=>X"00",
43699=>X"00",
43700=>X"00",
43701=>X"00",
43702=>X"00",
43703=>X"00",
43704=>X"00",
43705=>X"00",
43706=>X"00",
43707=>X"00",
43708=>X"00",
43709=>X"00",
43710=>X"00",
43711=>X"00",
43712=>X"00",
43713=>X"00",
43714=>X"00",
43715=>X"00",
43716=>X"00",
43717=>X"00",
43718=>X"00",
43719=>X"00",
43720=>X"00",
43721=>X"00",
43722=>X"00",
43723=>X"00",
43724=>X"00",
43725=>X"00",
43726=>X"00",
43727=>X"00",
43728=>X"00",
43729=>X"00",
43730=>X"00",
43731=>X"00",
43732=>X"00",
43733=>X"00",
43734=>X"00",
43735=>X"00",
43736=>X"00",
43737=>X"00",
43738=>X"00",
43739=>X"00",
43740=>X"00",
43741=>X"00",
43742=>X"00",
43743=>X"00",
43744=>X"00",
43745=>X"00",
43746=>X"00",
43747=>X"00",
43748=>X"00",
43749=>X"00",
43750=>X"00",
43751=>X"00",
43752=>X"00",
43753=>X"00",
43754=>X"00",
43755=>X"00",
43756=>X"00",
43757=>X"00",
43758=>X"00",
43759=>X"00",
43760=>X"00",
43761=>X"00",
43762=>X"00",
43763=>X"00",
43764=>X"00",
43765=>X"00",
43766=>X"00",
43767=>X"00",
43768=>X"00",
43769=>X"00",
43770=>X"00",
43771=>X"00",
43772=>X"00",
43773=>X"00",
43774=>X"00",
43775=>X"00",
43776=>X"00",
43777=>X"00",
43778=>X"00",
43779=>X"00",
43780=>X"00",
43781=>X"00",
43782=>X"00",
43783=>X"00",
43784=>X"00",
43785=>X"00",
43786=>X"00",
43787=>X"00",
43788=>X"00",
43789=>X"00",
43790=>X"00",
43791=>X"00",
43792=>X"00",
43793=>X"00",
43794=>X"00",
43795=>X"00",
43796=>X"00",
43797=>X"00",
43798=>X"00",
43799=>X"00",
43800=>X"00",
43801=>X"00",
43802=>X"00",
43803=>X"00",
43804=>X"00",
43805=>X"00",
43806=>X"00",
43807=>X"00",
43808=>X"00",
43809=>X"00",
43810=>X"00",
43811=>X"00",
43812=>X"00",
43813=>X"00",
43814=>X"00",
43815=>X"00",
43816=>X"00",
43817=>X"00",
43818=>X"00",
43819=>X"00",
43820=>X"00",
43821=>X"00",
43822=>X"00",
43823=>X"00",
43824=>X"00",
43825=>X"00",
43826=>X"00",
43827=>X"00",
43828=>X"00",
43829=>X"00",
43830=>X"00",
43831=>X"00",
43832=>X"00",
43833=>X"00",
43834=>X"00",
43835=>X"00",
43836=>X"00",
43837=>X"00",
43838=>X"00",
43839=>X"00",
43840=>X"00",
43841=>X"00",
43842=>X"00",
43843=>X"00",
43844=>X"00",
43845=>X"00",
43846=>X"00",
43847=>X"00",
43848=>X"00",
43849=>X"00",
43850=>X"00",
43851=>X"00",
43852=>X"00",
43853=>X"00",
43854=>X"00",
43855=>X"00",
43856=>X"00",
43857=>X"00",
43858=>X"00",
43859=>X"00",
43860=>X"00",
43861=>X"00",
43862=>X"00",
43863=>X"00",
43864=>X"00",
43865=>X"00",
43866=>X"00",
43867=>X"00",
43868=>X"00",
43869=>X"00",
43870=>X"00",
43871=>X"00",
43872=>X"00",
43873=>X"00",
43874=>X"00",
43875=>X"00",
43876=>X"00",
43877=>X"00",
43878=>X"00",
43879=>X"00",
43880=>X"00",
43881=>X"00",
43882=>X"00",
43883=>X"00",
43884=>X"00",
43885=>X"00",
43886=>X"00",
43887=>X"00",
43888=>X"00",
43889=>X"00",
43890=>X"00",
43891=>X"00",
43892=>X"00",
43893=>X"00",
43894=>X"00",
43895=>X"00",
43896=>X"00",
43897=>X"00",
43898=>X"00",
43899=>X"00",
43900=>X"00",
43901=>X"00",
43902=>X"00",
43903=>X"00",
43904=>X"00",
43905=>X"00",
43906=>X"00",
43907=>X"00",
43908=>X"00",
43909=>X"00",
43910=>X"00",
43911=>X"00",
43912=>X"00",
43913=>X"00",
43914=>X"00",
43915=>X"00",
43916=>X"00",
43917=>X"00",
43918=>X"00",
43919=>X"00",
43920=>X"00",
43921=>X"00",
43922=>X"00",
43923=>X"00",
43924=>X"00",
43925=>X"00",
43926=>X"00",
43927=>X"00",
43928=>X"00",
43929=>X"00",
43930=>X"00",
43931=>X"00",
43932=>X"00",
43933=>X"00",
43934=>X"00",
43935=>X"00",
43936=>X"00",
43937=>X"00",
43938=>X"00",
43939=>X"00",
43940=>X"00",
43941=>X"00",
43942=>X"00",
43943=>X"00",
43944=>X"00",
43945=>X"00",
43946=>X"00",
43947=>X"00",
43948=>X"00",
43949=>X"00",
43950=>X"00",
43951=>X"00",
43952=>X"00",
43953=>X"00",
43954=>X"00",
43955=>X"00",
43956=>X"00",
43957=>X"00",
43958=>X"00",
43959=>X"00",
43960=>X"00",
43961=>X"00",
43962=>X"00",
43963=>X"00",
43964=>X"00",
43965=>X"00",
43966=>X"00",
43967=>X"00",
43968=>X"00",
43969=>X"00",
43970=>X"00",
43971=>X"00",
43972=>X"00",
43973=>X"00",
43974=>X"00",
43975=>X"00",
43976=>X"00",
43977=>X"00",
43978=>X"00",
43979=>X"00",
43980=>X"00",
43981=>X"00",
43982=>X"00",
43983=>X"00",
43984=>X"00",
43985=>X"00",
43986=>X"00",
43987=>X"00",
43988=>X"00",
43989=>X"00",
43990=>X"00",
43991=>X"00",
43992=>X"00",
43993=>X"00",
43994=>X"00",
43995=>X"00",
43996=>X"00",
43997=>X"00",
43998=>X"00",
43999=>X"00",
44000=>X"00",
44001=>X"00",
44002=>X"00",
44003=>X"00",
44004=>X"00",
44005=>X"00",
44006=>X"00",
44007=>X"00",
44008=>X"00",
44009=>X"00",
44010=>X"00",
44011=>X"00",
44012=>X"00",
44013=>X"00",
44014=>X"00",
44015=>X"00",
44016=>X"00",
44017=>X"00",
44018=>X"00",
44019=>X"00",
44020=>X"00",
44021=>X"00",
44022=>X"00",
44023=>X"00",
44024=>X"00",
44025=>X"00",
44026=>X"00",
44027=>X"00",
44028=>X"00",
44029=>X"00",
44030=>X"00",
44031=>X"00",
44032=>X"00",
44033=>X"00",
44034=>X"00",
44035=>X"00",
44036=>X"00",
44037=>X"00",
44038=>X"00",
44039=>X"00",
44040=>X"00",
44041=>X"00",
44042=>X"00",
44043=>X"00",
44044=>X"00",
44045=>X"00",
44046=>X"00",
44047=>X"00",
44048=>X"00",
44049=>X"00",
44050=>X"00",
44051=>X"00",
44052=>X"00",
44053=>X"00",
44054=>X"00",
44055=>X"00",
44056=>X"00",
44057=>X"00",
44058=>X"00",
44059=>X"00",
44060=>X"00",
44061=>X"00",
44062=>X"00",
44063=>X"00",
44064=>X"00",
44065=>X"00",
44066=>X"00",
44067=>X"00",
44068=>X"00",
44069=>X"00",
44070=>X"00",
44071=>X"00",
44072=>X"00",
44073=>X"00",
44074=>X"00",
44075=>X"00",
44076=>X"00",
44077=>X"00",
44078=>X"00",
44079=>X"00",
44080=>X"00",
44081=>X"00",
44082=>X"00",
44083=>X"00",
44084=>X"00",
44085=>X"00",
44086=>X"00",
44087=>X"00",
44088=>X"00",
44089=>X"00",
44090=>X"00",
44091=>X"00",
44092=>X"00",
44093=>X"00",
44094=>X"00",
44095=>X"00",
44096=>X"00",
44097=>X"00",
44098=>X"00",
44099=>X"00",
44100=>X"00",
44101=>X"00",
44102=>X"00",
44103=>X"00",
44104=>X"00",
44105=>X"00",
44106=>X"00",
44107=>X"00",
44108=>X"00",
44109=>X"00",
44110=>X"00",
44111=>X"00",
44112=>X"00",
44113=>X"00",
44114=>X"00",
44115=>X"00",
44116=>X"00",
44117=>X"00",
44118=>X"00",
44119=>X"00",
44120=>X"00",
44121=>X"00",
44122=>X"00",
44123=>X"00",
44124=>X"00",
44125=>X"00",
44126=>X"00",
44127=>X"00",
44128=>X"00",
44129=>X"00",
44130=>X"00",
44131=>X"00",
44132=>X"00",
44133=>X"00",
44134=>X"00",
44135=>X"00",
44136=>X"00",
44137=>X"00",
44138=>X"00",
44139=>X"00",
44140=>X"00",
44141=>X"00",
44142=>X"00",
44143=>X"00",
44144=>X"00",
44145=>X"00",
44146=>X"00",
44147=>X"00",
44148=>X"00",
44149=>X"00",
44150=>X"00",
44151=>X"00",
44152=>X"00",
44153=>X"00",
44154=>X"00",
44155=>X"00",
44156=>X"00",
44157=>X"00",
44158=>X"00",
44159=>X"00",
44160=>X"00",
44161=>X"00",
44162=>X"00",
44163=>X"00",
44164=>X"00",
44165=>X"00",
44166=>X"00",
44167=>X"00",
44168=>X"00",
44169=>X"00",
44170=>X"00",
44171=>X"00",
44172=>X"00",
44173=>X"00",
44174=>X"00",
44175=>X"00",
44176=>X"00",
44177=>X"00",
44178=>X"00",
44179=>X"00",
44180=>X"00",
44181=>X"00",
44182=>X"00",
44183=>X"00",
44184=>X"00",
44185=>X"00",
44186=>X"00",
44187=>X"00",
44188=>X"00",
44189=>X"00",
44190=>X"00",
44191=>X"00",
44192=>X"00",
44193=>X"00",
44194=>X"00",
44195=>X"00",
44196=>X"00",
44197=>X"00",
44198=>X"00",
44199=>X"00",
44200=>X"00",
44201=>X"00",
44202=>X"00",
44203=>X"00",
44204=>X"00",
44205=>X"00",
44206=>X"00",
44207=>X"00",
44208=>X"00",
44209=>X"00",
44210=>X"00",
44211=>X"00",
44212=>X"00",
44213=>X"00",
44214=>X"00",
44215=>X"00",
44216=>X"00",
44217=>X"00",
44218=>X"00",
44219=>X"00",
44220=>X"00",
44221=>X"00",
44222=>X"00",
44223=>X"00",
44224=>X"00",
44225=>X"00",
44226=>X"00",
44227=>X"00",
44228=>X"00",
44229=>X"00",
44230=>X"00",
44231=>X"00",
44232=>X"00",
44233=>X"00",
44234=>X"00",
44235=>X"00",
44236=>X"00",
44237=>X"00",
44238=>X"00",
44239=>X"00",
44240=>X"00",
44241=>X"00",
44242=>X"00",
44243=>X"00",
44244=>X"00",
44245=>X"00",
44246=>X"00",
44247=>X"00",
44248=>X"00",
44249=>X"00",
44250=>X"00",
44251=>X"00",
44252=>X"00",
44253=>X"00",
44254=>X"00",
44255=>X"00",
44256=>X"00",
44257=>X"00",
44258=>X"00",
44259=>X"00",
44260=>X"00",
44261=>X"00",
44262=>X"00",
44263=>X"00",
44264=>X"00",
44265=>X"00",
44266=>X"00",
44267=>X"00",
44268=>X"00",
44269=>X"00",
44270=>X"00",
44271=>X"00",
44272=>X"00",
44273=>X"00",
44274=>X"00",
44275=>X"00",
44276=>X"00",
44277=>X"00",
44278=>X"00",
44279=>X"00",
44280=>X"00",
44281=>X"00",
44282=>X"00",
44283=>X"00",
44284=>X"00",
44285=>X"00",
44286=>X"00",
44287=>X"00",
44288=>X"00",
44289=>X"00",
44290=>X"00",
44291=>X"00",
44292=>X"00",
44293=>X"00",
44294=>X"00",
44295=>X"00",
44296=>X"00",
44297=>X"00",
44298=>X"00",
44299=>X"00",
44300=>X"00",
44301=>X"00",
44302=>X"00",
44303=>X"00",
44304=>X"00",
44305=>X"00",
44306=>X"00",
44307=>X"00",
44308=>X"00",
44309=>X"00",
44310=>X"00",
44311=>X"00",
44312=>X"00",
44313=>X"00",
44314=>X"00",
44315=>X"00",
44316=>X"00",
44317=>X"00",
44318=>X"00",
44319=>X"00",
44320=>X"00",
44321=>X"00",
44322=>X"00",
44323=>X"00",
44324=>X"00",
44325=>X"00",
44326=>X"00",
44327=>X"00",
44328=>X"00",
44329=>X"00",
44330=>X"00",
44331=>X"00",
44332=>X"00",
44333=>X"00",
44334=>X"00",
44335=>X"00",
44336=>X"00",
44337=>X"00",
44338=>X"00",
44339=>X"00",
44340=>X"00",
44341=>X"00",
44342=>X"00",
44343=>X"00",
44344=>X"00",
44345=>X"00",
44346=>X"00",
44347=>X"00",
44348=>X"00",
44349=>X"00",
44350=>X"00",
44351=>X"00",
44352=>X"00",
44353=>X"00",
44354=>X"00",
44355=>X"00",
44356=>X"00",
44357=>X"00",
44358=>X"00",
44359=>X"00",
44360=>X"00",
44361=>X"00",
44362=>X"00",
44363=>X"00",
44364=>X"00",
44365=>X"00",
44366=>X"00",
44367=>X"00",
44368=>X"00",
44369=>X"00",
44370=>X"00",
44371=>X"00",
44372=>X"00",
44373=>X"00",
44374=>X"00",
44375=>X"00",
44376=>X"00",
44377=>X"00",
44378=>X"00",
44379=>X"00",
44380=>X"00",
44381=>X"00",
44382=>X"00",
44383=>X"00",
44384=>X"00",
44385=>X"00",
44386=>X"00",
44387=>X"00",
44388=>X"00",
44389=>X"00",
44390=>X"00",
44391=>X"00",
44392=>X"00",
44393=>X"00",
44394=>X"00",
44395=>X"00",
44396=>X"00",
44397=>X"00",
44398=>X"00",
44399=>X"00",
44400=>X"00",
44401=>X"00",
44402=>X"00",
44403=>X"00",
44404=>X"00",
44405=>X"00",
44406=>X"00",
44407=>X"00",
44408=>X"00",
44409=>X"00",
44410=>X"00",
44411=>X"00",
44412=>X"00",
44413=>X"00",
44414=>X"00",
44415=>X"00",
44416=>X"00",
44417=>X"00",
44418=>X"00",
44419=>X"00",
44420=>X"00",
44421=>X"00",
44422=>X"00",
44423=>X"00",
44424=>X"00",
44425=>X"00",
44426=>X"00",
44427=>X"00",
44428=>X"00",
44429=>X"00",
44430=>X"00",
44431=>X"00",
44432=>X"00",
44433=>X"00",
44434=>X"00",
44435=>X"00",
44436=>X"00",
44437=>X"00",
44438=>X"00",
44439=>X"00",
44440=>X"00",
44441=>X"00",
44442=>X"00",
44443=>X"00",
44444=>X"00",
44445=>X"00",
44446=>X"00",
44447=>X"00",
44448=>X"00",
44449=>X"00",
44450=>X"00",
44451=>X"00",
44452=>X"00",
44453=>X"00",
44454=>X"00",
44455=>X"00",
44456=>X"00",
44457=>X"00",
44458=>X"00",
44459=>X"00",
44460=>X"00",
44461=>X"00",
44462=>X"00",
44463=>X"00",
44464=>X"00",
44465=>X"00",
44466=>X"00",
44467=>X"00",
44468=>X"00",
44469=>X"00",
44470=>X"00",
44471=>X"00",
44472=>X"00",
44473=>X"00",
44474=>X"00",
44475=>X"00",
44476=>X"00",
44477=>X"00",
44478=>X"00",
44479=>X"00",
44480=>X"00",
44481=>X"00",
44482=>X"00",
44483=>X"00",
44484=>X"00",
44485=>X"00",
44486=>X"00",
44487=>X"00",
44488=>X"00",
44489=>X"00",
44490=>X"00",
44491=>X"00",
44492=>X"00",
44493=>X"00",
44494=>X"00",
44495=>X"00",
44496=>X"00",
44497=>X"00",
44498=>X"00",
44499=>X"00",
44500=>X"00",
44501=>X"00",
44502=>X"00",
44503=>X"00",
44504=>X"00",
44505=>X"00",
44506=>X"00",
44507=>X"00",
44508=>X"00",
44509=>X"00",
44510=>X"00",
44511=>X"00",
44512=>X"00",
44513=>X"00",
44514=>X"00",
44515=>X"00",
44516=>X"00",
44517=>X"00",
44518=>X"00",
44519=>X"00",
44520=>X"00",
44521=>X"00",
44522=>X"00",
44523=>X"00",
44524=>X"00",
44525=>X"00",
44526=>X"00",
44527=>X"00",
44528=>X"00",
44529=>X"00",
44530=>X"00",
44531=>X"00",
44532=>X"00",
44533=>X"00",
44534=>X"00",
44535=>X"00",
44536=>X"00",
44537=>X"00",
44538=>X"00",
44539=>X"00",
44540=>X"00",
44541=>X"00",
44542=>X"00",
44543=>X"00",
44544=>X"00",
44545=>X"00",
44546=>X"00",
44547=>X"00",
44548=>X"00",
44549=>X"00",
44550=>X"00",
44551=>X"00",
44552=>X"00",
44553=>X"00",
44554=>X"00",
44555=>X"00",
44556=>X"00",
44557=>X"00",
44558=>X"00",
44559=>X"00",
44560=>X"00",
44561=>X"00",
44562=>X"00",
44563=>X"00",
44564=>X"00",
44565=>X"00",
44566=>X"00",
44567=>X"00",
44568=>X"00",
44569=>X"00",
44570=>X"00",
44571=>X"00",
44572=>X"00",
44573=>X"00",
44574=>X"00",
44575=>X"00",
44576=>X"00",
44577=>X"00",
44578=>X"00",
44579=>X"00",
44580=>X"00",
44581=>X"00",
44582=>X"00",
44583=>X"00",
44584=>X"00",
44585=>X"00",
44586=>X"00",
44587=>X"00",
44588=>X"00",
44589=>X"00",
44590=>X"00",
44591=>X"00",
44592=>X"00",
44593=>X"00",
44594=>X"00",
44595=>X"00",
44596=>X"00",
44597=>X"00",
44598=>X"00",
44599=>X"00",
44600=>X"00",
44601=>X"00",
44602=>X"00",
44603=>X"00",
44604=>X"00",
44605=>X"00",
44606=>X"00",
44607=>X"00",
44608=>X"00",
44609=>X"00",
44610=>X"00",
44611=>X"00",
44612=>X"00",
44613=>X"00",
44614=>X"00",
44615=>X"00",
44616=>X"00",
44617=>X"00",
44618=>X"00",
44619=>X"00",
44620=>X"00",
44621=>X"00",
44622=>X"00",
44623=>X"00",
44624=>X"00",
44625=>X"00",
44626=>X"00",
44627=>X"00",
44628=>X"00",
44629=>X"00",
44630=>X"00",
44631=>X"00",
44632=>X"00",
44633=>X"00",
44634=>X"00",
44635=>X"00",
44636=>X"00",
44637=>X"00",
44638=>X"00",
44639=>X"00",
44640=>X"00",
44641=>X"00",
44642=>X"00",
44643=>X"00",
44644=>X"00",
44645=>X"00",
44646=>X"00",
44647=>X"00",
44648=>X"00",
44649=>X"00",
44650=>X"00",
44651=>X"00",
44652=>X"00",
44653=>X"00",
44654=>X"00",
44655=>X"00",
44656=>X"00",
44657=>X"00",
44658=>X"00",
44659=>X"00",
44660=>X"00",
44661=>X"00",
44662=>X"00",
44663=>X"00",
44664=>X"00",
44665=>X"00",
44666=>X"00",
44667=>X"00",
44668=>X"00",
44669=>X"00",
44670=>X"00",
44671=>X"00",
44672=>X"00",
44673=>X"00",
44674=>X"00",
44675=>X"00",
44676=>X"00",
44677=>X"00",
44678=>X"00",
44679=>X"00",
44680=>X"00",
44681=>X"00",
44682=>X"00",
44683=>X"00",
44684=>X"00",
44685=>X"00",
44686=>X"00",
44687=>X"00",
44688=>X"00",
44689=>X"00",
44690=>X"00",
44691=>X"00",
44692=>X"00",
44693=>X"00",
44694=>X"00",
44695=>X"00",
44696=>X"00",
44697=>X"00",
44698=>X"00",
44699=>X"00",
44700=>X"00",
44701=>X"00",
44702=>X"00",
44703=>X"00",
44704=>X"00",
44705=>X"00",
44706=>X"00",
44707=>X"00",
44708=>X"00",
44709=>X"00",
44710=>X"00",
44711=>X"00",
44712=>X"00",
44713=>X"00",
44714=>X"00",
44715=>X"00",
44716=>X"00",
44717=>X"00",
44718=>X"00",
44719=>X"00",
44720=>X"00",
44721=>X"00",
44722=>X"00",
44723=>X"00",
44724=>X"00",
44725=>X"00",
44726=>X"00",
44727=>X"00",
44728=>X"00",
44729=>X"00",
44730=>X"00",
44731=>X"00",
44732=>X"00",
44733=>X"00",
44734=>X"00",
44735=>X"00",
44736=>X"00",
44737=>X"00",
44738=>X"00",
44739=>X"00",
44740=>X"00",
44741=>X"00",
44742=>X"00",
44743=>X"00",
44744=>X"00",
44745=>X"00",
44746=>X"00",
44747=>X"00",
44748=>X"00",
44749=>X"00",
44750=>X"00",
44751=>X"00",
44752=>X"00",
44753=>X"00",
44754=>X"00",
44755=>X"00",
44756=>X"00",
44757=>X"00",
44758=>X"00",
44759=>X"00",
44760=>X"00",
44761=>X"00",
44762=>X"00",
44763=>X"00",
44764=>X"00",
44765=>X"00",
44766=>X"00",
44767=>X"00",
44768=>X"00",
44769=>X"00",
44770=>X"00",
44771=>X"00",
44772=>X"00",
44773=>X"00",
44774=>X"00",
44775=>X"00",
44776=>X"00",
44777=>X"00",
44778=>X"00",
44779=>X"00",
44780=>X"00",
44781=>X"00",
44782=>X"00",
44783=>X"00",
44784=>X"00",
44785=>X"00",
44786=>X"00",
44787=>X"00",
44788=>X"00",
44789=>X"00",
44790=>X"00",
44791=>X"00",
44792=>X"00",
44793=>X"00",
44794=>X"00",
44795=>X"00",
44796=>X"00",
44797=>X"00",
44798=>X"00",
44799=>X"00",
44800=>X"00",
44801=>X"00",
44802=>X"00",
44803=>X"00",
44804=>X"00",
44805=>X"00",
44806=>X"00",
44807=>X"00",
44808=>X"00",
44809=>X"00",
44810=>X"00",
44811=>X"00",
44812=>X"00",
44813=>X"00",
44814=>X"00",
44815=>X"00",
44816=>X"00",
44817=>X"00",
44818=>X"00",
44819=>X"00",
44820=>X"00",
44821=>X"00",
44822=>X"00",
44823=>X"00",
44824=>X"00",
44825=>X"00",
44826=>X"00",
44827=>X"00",
44828=>X"00",
44829=>X"00",
44830=>X"00",
44831=>X"00",
44832=>X"00",
44833=>X"00",
44834=>X"00",
44835=>X"00",
44836=>X"00",
44837=>X"00",
44838=>X"00",
44839=>X"00",
44840=>X"00",
44841=>X"00",
44842=>X"00",
44843=>X"00",
44844=>X"00",
44845=>X"00",
44846=>X"00",
44847=>X"00",
44848=>X"00",
44849=>X"00",
44850=>X"00",
44851=>X"00",
44852=>X"00",
44853=>X"00",
44854=>X"00",
44855=>X"00",
44856=>X"00",
44857=>X"00",
44858=>X"00",
44859=>X"00",
44860=>X"00",
44861=>X"00",
44862=>X"00",
44863=>X"00",
44864=>X"00",
44865=>X"00",
44866=>X"00",
44867=>X"00",
44868=>X"00",
44869=>X"00",
44870=>X"00",
44871=>X"00",
44872=>X"00",
44873=>X"00",
44874=>X"00",
44875=>X"00",
44876=>X"00",
44877=>X"00",
44878=>X"00",
44879=>X"00",
44880=>X"00",
44881=>X"00",
44882=>X"00",
44883=>X"00",
44884=>X"00",
44885=>X"00",
44886=>X"00",
44887=>X"00",
44888=>X"00",
44889=>X"00",
44890=>X"00",
44891=>X"00",
44892=>X"00",
44893=>X"00",
44894=>X"00",
44895=>X"00",
44896=>X"00",
44897=>X"00",
44898=>X"00",
44899=>X"00",
44900=>X"00",
44901=>X"00",
44902=>X"00",
44903=>X"00",
44904=>X"00",
44905=>X"00",
44906=>X"00",
44907=>X"00",
44908=>X"00",
44909=>X"00",
44910=>X"00",
44911=>X"00",
44912=>X"00",
44913=>X"00",
44914=>X"00",
44915=>X"00",
44916=>X"00",
44917=>X"00",
44918=>X"00",
44919=>X"00",
44920=>X"00",
44921=>X"00",
44922=>X"00",
44923=>X"00",
44924=>X"00",
44925=>X"00",
44926=>X"00",
44927=>X"00",
44928=>X"00",
44929=>X"00",
44930=>X"00",
44931=>X"00",
44932=>X"00",
44933=>X"00",
44934=>X"00",
44935=>X"00",
44936=>X"00",
44937=>X"00",
44938=>X"00",
44939=>X"00",
44940=>X"00",
44941=>X"00",
44942=>X"00",
44943=>X"00",
44944=>X"00",
44945=>X"00",
44946=>X"00",
44947=>X"00",
44948=>X"00",
44949=>X"00",
44950=>X"00",
44951=>X"00",
44952=>X"00",
44953=>X"00",
44954=>X"00",
44955=>X"00",
44956=>X"00",
44957=>X"00",
44958=>X"00",
44959=>X"00",
44960=>X"00",
44961=>X"00",
44962=>X"00",
44963=>X"00",
44964=>X"00",
44965=>X"00",
44966=>X"00",
44967=>X"00",
44968=>X"00",
44969=>X"00",
44970=>X"00",
44971=>X"00",
44972=>X"00",
44973=>X"00",
44974=>X"00",
44975=>X"00",
44976=>X"00",
44977=>X"00",
44978=>X"00",
44979=>X"00",
44980=>X"00",
44981=>X"00",
44982=>X"00",
44983=>X"00",
44984=>X"00",
44985=>X"00",
44986=>X"00",
44987=>X"00",
44988=>X"00",
44989=>X"00",
44990=>X"00",
44991=>X"00",
44992=>X"00",
44993=>X"00",
44994=>X"00",
44995=>X"00",
44996=>X"00",
44997=>X"00",
44998=>X"00",
44999=>X"00",
45000=>X"00",
45001=>X"00",
45002=>X"00",
45003=>X"00",
45004=>X"00",
45005=>X"00",
45006=>X"00",
45007=>X"00",
45008=>X"00",
45009=>X"00",
45010=>X"00",
45011=>X"00",
45012=>X"00",
45013=>X"00",
45014=>X"00",
45015=>X"00",
45016=>X"00",
45017=>X"00",
45018=>X"00",
45019=>X"00",
45020=>X"00",
45021=>X"00",
45022=>X"00",
45023=>X"00",
45024=>X"00",
45025=>X"00",
45026=>X"00",
45027=>X"00",
45028=>X"00",
45029=>X"00",
45030=>X"00",
45031=>X"00",
45032=>X"00",
45033=>X"00",
45034=>X"00",
45035=>X"00",
45036=>X"00",
45037=>X"00",
45038=>X"00",
45039=>X"00",
45040=>X"00",
45041=>X"00",
45042=>X"00",
45043=>X"00",
45044=>X"00",
45045=>X"00",
45046=>X"00",
45047=>X"00",
45048=>X"00",
45049=>X"00",
45050=>X"00",
45051=>X"00",
45052=>X"00",
45053=>X"00",
45054=>X"00",
45055=>X"00",
45056=>X"00",
45057=>X"00",
45058=>X"00",
45059=>X"00",
45060=>X"00",
45061=>X"00",
45062=>X"00",
45063=>X"00",
45064=>X"00",
45065=>X"00",
45066=>X"00",
45067=>X"00",
45068=>X"00",
45069=>X"00",
45070=>X"00",
45071=>X"00",
45072=>X"00",
45073=>X"00",
45074=>X"00",
45075=>X"00",
45076=>X"00",
45077=>X"00",
45078=>X"00",
45079=>X"00",
45080=>X"00",
45081=>X"00",
45082=>X"00",
45083=>X"00",
45084=>X"00",
45085=>X"00",
45086=>X"00",
45087=>X"00",
45088=>X"00",
45089=>X"00",
45090=>X"00",
45091=>X"00",
45092=>X"00",
45093=>X"00",
45094=>X"00",
45095=>X"00",
45096=>X"00",
45097=>X"00",
45098=>X"00",
45099=>X"00",
45100=>X"00",
45101=>X"00",
45102=>X"00",
45103=>X"00",
45104=>X"00",
45105=>X"00",
45106=>X"00",
45107=>X"00",
45108=>X"00",
45109=>X"00",
45110=>X"00",
45111=>X"00",
45112=>X"00",
45113=>X"00",
45114=>X"00",
45115=>X"00",
45116=>X"00",
45117=>X"00",
45118=>X"00",
45119=>X"00",
45120=>X"00",
45121=>X"00",
45122=>X"00",
45123=>X"00",
45124=>X"00",
45125=>X"00",
45126=>X"00",
45127=>X"00",
45128=>X"00",
45129=>X"00",
45130=>X"00",
45131=>X"00",
45132=>X"00",
45133=>X"00",
45134=>X"00",
45135=>X"00",
45136=>X"00",
45137=>X"00",
45138=>X"00",
45139=>X"00",
45140=>X"00",
45141=>X"00",
45142=>X"00",
45143=>X"00",
45144=>X"00",
45145=>X"00",
45146=>X"00",
45147=>X"00",
45148=>X"00",
45149=>X"00",
45150=>X"00",
45151=>X"00",
45152=>X"00",
45153=>X"00",
45154=>X"00",
45155=>X"00",
45156=>X"00",
45157=>X"00",
45158=>X"00",
45159=>X"00",
45160=>X"00",
45161=>X"00",
45162=>X"00",
45163=>X"00",
45164=>X"00",
45165=>X"00",
45166=>X"00",
45167=>X"00",
45168=>X"00",
45169=>X"00",
45170=>X"00",
45171=>X"00",
45172=>X"00",
45173=>X"00",
45174=>X"00",
45175=>X"00",
45176=>X"00",
45177=>X"00",
45178=>X"00",
45179=>X"00",
45180=>X"00",
45181=>X"00",
45182=>X"00",
45183=>X"00",
45184=>X"00",
45185=>X"00",
45186=>X"00",
45187=>X"00",
45188=>X"00",
45189=>X"00",
45190=>X"00",
45191=>X"00",
45192=>X"00",
45193=>X"00",
45194=>X"00",
45195=>X"00",
45196=>X"00",
45197=>X"00",
45198=>X"00",
45199=>X"00",
45200=>X"00",
45201=>X"00",
45202=>X"00",
45203=>X"00",
45204=>X"00",
45205=>X"00",
45206=>X"00",
45207=>X"00",
45208=>X"00",
45209=>X"00",
45210=>X"00",
45211=>X"00",
45212=>X"00",
45213=>X"00",
45214=>X"00",
45215=>X"00",
45216=>X"00",
45217=>X"00",
45218=>X"00",
45219=>X"00",
45220=>X"00",
45221=>X"00",
45222=>X"00",
45223=>X"00",
45224=>X"00",
45225=>X"00",
45226=>X"00",
45227=>X"00",
45228=>X"00",
45229=>X"00",
45230=>X"00",
45231=>X"00",
45232=>X"00",
45233=>X"00",
45234=>X"00",
45235=>X"00",
45236=>X"00",
45237=>X"00",
45238=>X"00",
45239=>X"00",
45240=>X"00",
45241=>X"00",
45242=>X"00",
45243=>X"00",
45244=>X"00",
45245=>X"00",
45246=>X"00",
45247=>X"00",
45248=>X"00",
45249=>X"00",
45250=>X"00",
45251=>X"00",
45252=>X"00",
45253=>X"00",
45254=>X"00",
45255=>X"00",
45256=>X"00",
45257=>X"00",
45258=>X"00",
45259=>X"00",
45260=>X"00",
45261=>X"00",
45262=>X"00",
45263=>X"00",
45264=>X"00",
45265=>X"00",
45266=>X"00",
45267=>X"00",
45268=>X"00",
45269=>X"00",
45270=>X"00",
45271=>X"00",
45272=>X"00",
45273=>X"00",
45274=>X"00",
45275=>X"00",
45276=>X"00",
45277=>X"00",
45278=>X"00",
45279=>X"00",
45280=>X"00",
45281=>X"00",
45282=>X"00",
45283=>X"00",
45284=>X"00",
45285=>X"00",
45286=>X"00",
45287=>X"00",
45288=>X"00",
45289=>X"00",
45290=>X"00",
45291=>X"00",
45292=>X"00",
45293=>X"00",
45294=>X"00",
45295=>X"00",
45296=>X"00",
45297=>X"00",
45298=>X"00",
45299=>X"00",
45300=>X"00",
45301=>X"00",
45302=>X"00",
45303=>X"00",
45304=>X"00",
45305=>X"00",
45306=>X"00",
45307=>X"00",
45308=>X"00",
45309=>X"00",
45310=>X"00",
45311=>X"00",
45312=>X"00",
45313=>X"00",
45314=>X"00",
45315=>X"00",
45316=>X"00",
45317=>X"00",
45318=>X"00",
45319=>X"00",
45320=>X"00",
45321=>X"00",
45322=>X"00",
45323=>X"00",
45324=>X"00",
45325=>X"00",
45326=>X"00",
45327=>X"00",
45328=>X"00",
45329=>X"00",
45330=>X"00",
45331=>X"00",
45332=>X"00",
45333=>X"00",
45334=>X"00",
45335=>X"00",
45336=>X"00",
45337=>X"00",
45338=>X"00",
45339=>X"00",
45340=>X"00",
45341=>X"00",
45342=>X"00",
45343=>X"00",
45344=>X"00",
45345=>X"00",
45346=>X"00",
45347=>X"00",
45348=>X"00",
45349=>X"00",
45350=>X"00",
45351=>X"00",
45352=>X"00",
45353=>X"00",
45354=>X"00",
45355=>X"00",
45356=>X"00",
45357=>X"00",
45358=>X"00",
45359=>X"00",
45360=>X"00",
45361=>X"00",
45362=>X"00",
45363=>X"00",
45364=>X"00",
45365=>X"00",
45366=>X"00",
45367=>X"00",
45368=>X"00",
45369=>X"00",
45370=>X"00",
45371=>X"00",
45372=>X"00",
45373=>X"00",
45374=>X"00",
45375=>X"00",
45376=>X"00",
45377=>X"00",
45378=>X"00",
45379=>X"00",
45380=>X"00",
45381=>X"00",
45382=>X"00",
45383=>X"00",
45384=>X"00",
45385=>X"00",
45386=>X"00",
45387=>X"00",
45388=>X"00",
45389=>X"00",
45390=>X"00",
45391=>X"00",
45392=>X"00",
45393=>X"00",
45394=>X"00",
45395=>X"00",
45396=>X"00",
45397=>X"00",
45398=>X"00",
45399=>X"00",
45400=>X"00",
45401=>X"00",
45402=>X"00",
45403=>X"00",
45404=>X"00",
45405=>X"00",
45406=>X"00",
45407=>X"00",
45408=>X"00",
45409=>X"00",
45410=>X"00",
45411=>X"00",
45412=>X"00",
45413=>X"00",
45414=>X"00",
45415=>X"00",
45416=>X"00",
45417=>X"00",
45418=>X"00",
45419=>X"00",
45420=>X"00",
45421=>X"00",
45422=>X"00",
45423=>X"00",
45424=>X"00",
45425=>X"00",
45426=>X"00",
45427=>X"00",
45428=>X"00",
45429=>X"00",
45430=>X"00",
45431=>X"00",
45432=>X"00",
45433=>X"00",
45434=>X"00",
45435=>X"00",
45436=>X"00",
45437=>X"00",
45438=>X"00",
45439=>X"00",
45440=>X"00",
45441=>X"00",
45442=>X"00",
45443=>X"00",
45444=>X"00",
45445=>X"00",
45446=>X"00",
45447=>X"00",
45448=>X"00",
45449=>X"00",
45450=>X"00",
45451=>X"00",
45452=>X"00",
45453=>X"00",
45454=>X"00",
45455=>X"00",
45456=>X"00",
45457=>X"00",
45458=>X"00",
45459=>X"00",
45460=>X"00",
45461=>X"00",
45462=>X"00",
45463=>X"00",
45464=>X"00",
45465=>X"00",
45466=>X"00",
45467=>X"00",
45468=>X"00",
45469=>X"00",
45470=>X"00",
45471=>X"00",
45472=>X"00",
45473=>X"00",
45474=>X"00",
45475=>X"00",
45476=>X"00",
45477=>X"00",
45478=>X"00",
45479=>X"00",
45480=>X"00",
45481=>X"00",
45482=>X"00",
45483=>X"00",
45484=>X"00",
45485=>X"00",
45486=>X"00",
45487=>X"00",
45488=>X"00",
45489=>X"00",
45490=>X"00",
45491=>X"00",
45492=>X"00",
45493=>X"00",
45494=>X"00",
45495=>X"00",
45496=>X"00",
45497=>X"00",
45498=>X"00",
45499=>X"00",
45500=>X"00",
45501=>X"00",
45502=>X"00",
45503=>X"00",
45504=>X"00",
45505=>X"00",
45506=>X"00",
45507=>X"00",
45508=>X"00",
45509=>X"00",
45510=>X"00",
45511=>X"00",
45512=>X"00",
45513=>X"00",
45514=>X"00",
45515=>X"00",
45516=>X"00",
45517=>X"00",
45518=>X"00",
45519=>X"00",
45520=>X"00",
45521=>X"00",
45522=>X"00",
45523=>X"00",
45524=>X"00",
45525=>X"00",
45526=>X"00",
45527=>X"00",
45528=>X"00",
45529=>X"00",
45530=>X"00",
45531=>X"00",
45532=>X"00",
45533=>X"00",
45534=>X"00",
45535=>X"00",
45536=>X"00",
45537=>X"00",
45538=>X"00",
45539=>X"00",
45540=>X"00",
45541=>X"00",
45542=>X"00",
45543=>X"00",
45544=>X"00",
45545=>X"00",
45546=>X"00",
45547=>X"00",
45548=>X"00",
45549=>X"00",
45550=>X"00",
45551=>X"00",
45552=>X"00",
45553=>X"00",
45554=>X"00",
45555=>X"00",
45556=>X"00",
45557=>X"00",
45558=>X"00",
45559=>X"00",
45560=>X"00",
45561=>X"00",
45562=>X"00",
45563=>X"00",
45564=>X"00",
45565=>X"00",
45566=>X"00",
45567=>X"00",
45568=>X"00",
45569=>X"00",
45570=>X"00",
45571=>X"00",
45572=>X"00",
45573=>X"00",
45574=>X"00",
45575=>X"00",
45576=>X"00",
45577=>X"00",
45578=>X"00",
45579=>X"00",
45580=>X"00",
45581=>X"00",
45582=>X"00",
45583=>X"00",
45584=>X"00",
45585=>X"00",
45586=>X"00",
45587=>X"00",
45588=>X"00",
45589=>X"00",
45590=>X"00",
45591=>X"00",
45592=>X"00",
45593=>X"00",
45594=>X"00",
45595=>X"00",
45596=>X"00",
45597=>X"00",
45598=>X"00",
45599=>X"00",
45600=>X"00",
45601=>X"00",
45602=>X"00",
45603=>X"00",
45604=>X"00",
45605=>X"00",
45606=>X"00",
45607=>X"00",
45608=>X"00",
45609=>X"00",
45610=>X"00",
45611=>X"00",
45612=>X"00",
45613=>X"00",
45614=>X"00",
45615=>X"00",
45616=>X"00",
45617=>X"00",
45618=>X"00",
45619=>X"00",
45620=>X"00",
45621=>X"00",
45622=>X"00",
45623=>X"00",
45624=>X"00",
45625=>X"00",
45626=>X"00",
45627=>X"00",
45628=>X"00",
45629=>X"00",
45630=>X"00",
45631=>X"00",
45632=>X"00",
45633=>X"00",
45634=>X"00",
45635=>X"00",
45636=>X"00",
45637=>X"00",
45638=>X"00",
45639=>X"00",
45640=>X"00",
45641=>X"00",
45642=>X"00",
45643=>X"00",
45644=>X"00",
45645=>X"00",
45646=>X"00",
45647=>X"00",
45648=>X"00",
45649=>X"00",
45650=>X"00",
45651=>X"00",
45652=>X"00",
45653=>X"00",
45654=>X"00",
45655=>X"00",
45656=>X"00",
45657=>X"00",
45658=>X"00",
45659=>X"00",
45660=>X"00",
45661=>X"00",
45662=>X"00",
45663=>X"00",
45664=>X"00",
45665=>X"00",
45666=>X"00",
45667=>X"00",
45668=>X"00",
45669=>X"00",
45670=>X"00",
45671=>X"00",
45672=>X"00",
45673=>X"00",
45674=>X"00",
45675=>X"00",
45676=>X"00",
45677=>X"00",
45678=>X"00",
45679=>X"00",
45680=>X"00",
45681=>X"00",
45682=>X"00",
45683=>X"00",
45684=>X"00",
45685=>X"00",
45686=>X"00",
45687=>X"00",
45688=>X"00",
45689=>X"00",
45690=>X"00",
45691=>X"00",
45692=>X"00",
45693=>X"00",
45694=>X"00",
45695=>X"00",
45696=>X"00",
45697=>X"00",
45698=>X"00",
45699=>X"00",
45700=>X"00",
45701=>X"00",
45702=>X"00",
45703=>X"00",
45704=>X"00",
45705=>X"00",
45706=>X"00",
45707=>X"00",
45708=>X"00",
45709=>X"00",
45710=>X"00",
45711=>X"00",
45712=>X"00",
45713=>X"00",
45714=>X"00",
45715=>X"00",
45716=>X"00",
45717=>X"00",
45718=>X"00",
45719=>X"00",
45720=>X"00",
45721=>X"00",
45722=>X"00",
45723=>X"00",
45724=>X"00",
45725=>X"00",
45726=>X"00",
45727=>X"00",
45728=>X"00",
45729=>X"00",
45730=>X"00",
45731=>X"00",
45732=>X"00",
45733=>X"00",
45734=>X"00",
45735=>X"00",
45736=>X"00",
45737=>X"00",
45738=>X"00",
45739=>X"00",
45740=>X"00",
45741=>X"00",
45742=>X"00",
45743=>X"00",
45744=>X"00",
45745=>X"00",
45746=>X"00",
45747=>X"00",
45748=>X"00",
45749=>X"00",
45750=>X"00",
45751=>X"00",
45752=>X"00",
45753=>X"00",
45754=>X"00",
45755=>X"00",
45756=>X"00",
45757=>X"00",
45758=>X"00",
45759=>X"00",
45760=>X"00",
45761=>X"00",
45762=>X"00",
45763=>X"00",
45764=>X"00",
45765=>X"00",
45766=>X"00",
45767=>X"00",
45768=>X"00",
45769=>X"00",
45770=>X"00",
45771=>X"00",
45772=>X"00",
45773=>X"00",
45774=>X"00",
45775=>X"00",
45776=>X"00",
45777=>X"00",
45778=>X"00",
45779=>X"00",
45780=>X"00",
45781=>X"00",
45782=>X"00",
45783=>X"00",
45784=>X"00",
45785=>X"00",
45786=>X"00",
45787=>X"00",
45788=>X"00",
45789=>X"00",
45790=>X"00",
45791=>X"00",
45792=>X"00",
45793=>X"00",
45794=>X"00",
45795=>X"00",
45796=>X"00",
45797=>X"00",
45798=>X"00",
45799=>X"00",
45800=>X"00",
45801=>X"00",
45802=>X"00",
45803=>X"00",
45804=>X"00",
45805=>X"00",
45806=>X"00",
45807=>X"00",
45808=>X"00",
45809=>X"00",
45810=>X"00",
45811=>X"00",
45812=>X"00",
45813=>X"00",
45814=>X"00",
45815=>X"00",
45816=>X"00",
45817=>X"00",
45818=>X"00",
45819=>X"00",
45820=>X"00",
45821=>X"00",
45822=>X"00",
45823=>X"00",
45824=>X"00",
45825=>X"00",
45826=>X"00",
45827=>X"00",
45828=>X"00",
45829=>X"00",
45830=>X"00",
45831=>X"00",
45832=>X"00",
45833=>X"00",
45834=>X"00",
45835=>X"00",
45836=>X"00",
45837=>X"00",
45838=>X"00",
45839=>X"00",
45840=>X"00",
45841=>X"00",
45842=>X"00",
45843=>X"00",
45844=>X"00",
45845=>X"00",
45846=>X"00",
45847=>X"00",
45848=>X"00",
45849=>X"00",
45850=>X"00",
45851=>X"00",
45852=>X"00",
45853=>X"00",
45854=>X"00",
45855=>X"00",
45856=>X"00",
45857=>X"00",
45858=>X"00",
45859=>X"00",
45860=>X"00",
45861=>X"00",
45862=>X"00",
45863=>X"00",
45864=>X"00",
45865=>X"00",
45866=>X"00",
45867=>X"00",
45868=>X"00",
45869=>X"00",
45870=>X"00",
45871=>X"00",
45872=>X"00",
45873=>X"00",
45874=>X"00",
45875=>X"00",
45876=>X"00",
45877=>X"00",
45878=>X"00",
45879=>X"00",
45880=>X"00",
45881=>X"00",
45882=>X"00",
45883=>X"00",
45884=>X"00",
45885=>X"00",
45886=>X"00",
45887=>X"00",
45888=>X"00",
45889=>X"00",
45890=>X"00",
45891=>X"00",
45892=>X"00",
45893=>X"00",
45894=>X"00",
45895=>X"00",
45896=>X"00",
45897=>X"00",
45898=>X"00",
45899=>X"00",
45900=>X"00",
45901=>X"00",
45902=>X"00",
45903=>X"00",
45904=>X"00",
45905=>X"00",
45906=>X"00",
45907=>X"00",
45908=>X"00",
45909=>X"00",
45910=>X"00",
45911=>X"00",
45912=>X"00",
45913=>X"00",
45914=>X"00",
45915=>X"00",
45916=>X"00",
45917=>X"00",
45918=>X"00",
45919=>X"00",
45920=>X"00",
45921=>X"00",
45922=>X"00",
45923=>X"00",
45924=>X"00",
45925=>X"00",
45926=>X"00",
45927=>X"00",
45928=>X"00",
45929=>X"00",
45930=>X"00",
45931=>X"00",
45932=>X"00",
45933=>X"00",
45934=>X"00",
45935=>X"00",
45936=>X"00",
45937=>X"00",
45938=>X"00",
45939=>X"00",
45940=>X"00",
45941=>X"00",
45942=>X"00",
45943=>X"00",
45944=>X"00",
45945=>X"00",
45946=>X"00",
45947=>X"00",
45948=>X"00",
45949=>X"00",
45950=>X"00",
45951=>X"00",
45952=>X"00",
45953=>X"00",
45954=>X"00",
45955=>X"00",
45956=>X"00",
45957=>X"00",
45958=>X"00",
45959=>X"00",
45960=>X"00",
45961=>X"00",
45962=>X"00",
45963=>X"00",
45964=>X"00",
45965=>X"00",
45966=>X"00",
45967=>X"00",
45968=>X"00",
45969=>X"00",
45970=>X"00",
45971=>X"00",
45972=>X"00",
45973=>X"00",
45974=>X"00",
45975=>X"00",
45976=>X"00",
45977=>X"00",
45978=>X"00",
45979=>X"00",
45980=>X"00",
45981=>X"00",
45982=>X"00",
45983=>X"00",
45984=>X"00",
45985=>X"00",
45986=>X"00",
45987=>X"00",
45988=>X"00",
45989=>X"00",
45990=>X"00",
45991=>X"00",
45992=>X"00",
45993=>X"00",
45994=>X"00",
45995=>X"00",
45996=>X"00",
45997=>X"00",
45998=>X"00",
45999=>X"00",
46000=>X"00",
46001=>X"00",
46002=>X"00",
46003=>X"00",
46004=>X"00",
46005=>X"00",
46006=>X"00",
46007=>X"00",
46008=>X"00",
46009=>X"00",
46010=>X"00",
46011=>X"00",
46012=>X"00",
46013=>X"00",
46014=>X"00",
46015=>X"00",
46016=>X"00",
46017=>X"00",
46018=>X"00",
46019=>X"00",
46020=>X"00",
46021=>X"00",
46022=>X"00",
46023=>X"00",
46024=>X"00",
46025=>X"00",
46026=>X"00",
46027=>X"00",
46028=>X"00",
46029=>X"00",
46030=>X"00",
46031=>X"00",
46032=>X"00",
46033=>X"00",
46034=>X"00",
46035=>X"00",
46036=>X"00",
46037=>X"00",
46038=>X"00",
46039=>X"00",
46040=>X"00",
46041=>X"00",
46042=>X"00",
46043=>X"00",
46044=>X"00",
46045=>X"00",
46046=>X"00",
46047=>X"00",
46048=>X"00",
46049=>X"00",
46050=>X"00",
46051=>X"00",
46052=>X"00",
46053=>X"00",
46054=>X"00",
46055=>X"00",
46056=>X"00",
46057=>X"00",
46058=>X"00",
46059=>X"00",
46060=>X"00",
46061=>X"00",
46062=>X"00",
46063=>X"00",
46064=>X"00",
46065=>X"00",
46066=>X"00",
46067=>X"00",
46068=>X"00",
46069=>X"00",
46070=>X"00",
46071=>X"00",
46072=>X"00",
46073=>X"00",
46074=>X"00",
46075=>X"00",
46076=>X"00",
46077=>X"00",
46078=>X"00",
46079=>X"00",
46080=>X"00",
46081=>X"00",
46082=>X"00",
46083=>X"00",
46084=>X"00",
46085=>X"00",
46086=>X"00",
46087=>X"00",
46088=>X"00",
46089=>X"00",
46090=>X"00",
46091=>X"00",
46092=>X"00",
46093=>X"00",
46094=>X"00",
46095=>X"00",
46096=>X"00",
46097=>X"00",
46098=>X"00",
46099=>X"00",
46100=>X"00",
46101=>X"00",
46102=>X"00",
46103=>X"00",
46104=>X"00",
46105=>X"00",
46106=>X"00",
46107=>X"00",
46108=>X"00",
46109=>X"00",
46110=>X"00",
46111=>X"00",
46112=>X"00",
46113=>X"00",
46114=>X"00",
46115=>X"00",
46116=>X"00",
46117=>X"00",
46118=>X"00",
46119=>X"00",
46120=>X"00",
46121=>X"00",
46122=>X"00",
46123=>X"00",
46124=>X"00",
46125=>X"00",
46126=>X"00",
46127=>X"00",
46128=>X"00",
46129=>X"00",
46130=>X"00",
46131=>X"00",
46132=>X"00",
46133=>X"00",
46134=>X"00",
46135=>X"00",
46136=>X"00",
46137=>X"00",
46138=>X"00",
46139=>X"00",
46140=>X"00",
46141=>X"00",
46142=>X"00",
46143=>X"00",
46144=>X"00",
46145=>X"00",
46146=>X"00",
46147=>X"00",
46148=>X"00",
46149=>X"00",
46150=>X"00",
46151=>X"00",
46152=>X"00",
46153=>X"00",
46154=>X"00",
46155=>X"00",
46156=>X"00",
46157=>X"00",
46158=>X"00",
46159=>X"00",
46160=>X"00",
46161=>X"00",
46162=>X"00",
46163=>X"00",
46164=>X"00",
46165=>X"00",
46166=>X"00",
46167=>X"00",
46168=>X"00",
46169=>X"00",
46170=>X"00",
46171=>X"00",
46172=>X"00",
46173=>X"00",
46174=>X"00",
46175=>X"00",
46176=>X"00",
46177=>X"00",
46178=>X"00",
46179=>X"00",
46180=>X"00",
46181=>X"00",
46182=>X"00",
46183=>X"00",
46184=>X"00",
46185=>X"00",
46186=>X"00",
46187=>X"00",
46188=>X"00",
46189=>X"00",
46190=>X"00",
46191=>X"00",
46192=>X"00",
46193=>X"00",
46194=>X"00",
46195=>X"00",
46196=>X"00",
46197=>X"00",
46198=>X"00",
46199=>X"00",
46200=>X"00",
46201=>X"00",
46202=>X"00",
46203=>X"00",
46204=>X"00",
46205=>X"00",
46206=>X"00",
46207=>X"00",
46208=>X"00",
46209=>X"00",
46210=>X"00",
46211=>X"00",
46212=>X"00",
46213=>X"00",
46214=>X"00",
46215=>X"00",
46216=>X"00",
46217=>X"00",
46218=>X"00",
46219=>X"00",
46220=>X"00",
46221=>X"00",
46222=>X"00",
46223=>X"00",
46224=>X"00",
46225=>X"00",
46226=>X"00",
46227=>X"00",
46228=>X"00",
46229=>X"00",
46230=>X"00",
46231=>X"00",
46232=>X"00",
46233=>X"00",
46234=>X"00",
46235=>X"00",
46236=>X"00",
46237=>X"00",
46238=>X"00",
46239=>X"00",
46240=>X"00",
46241=>X"00",
46242=>X"00",
46243=>X"00",
46244=>X"00",
46245=>X"00",
46246=>X"00",
46247=>X"00",
46248=>X"00",
46249=>X"00",
46250=>X"00",
46251=>X"00",
46252=>X"00",
46253=>X"00",
46254=>X"00",
46255=>X"00",
46256=>X"00",
46257=>X"00",
46258=>X"00",
46259=>X"00",
46260=>X"00",
46261=>X"00",
46262=>X"00",
46263=>X"00",
46264=>X"00",
46265=>X"00",
46266=>X"00",
46267=>X"00",
46268=>X"00",
46269=>X"00",
46270=>X"00",
46271=>X"00",
46272=>X"00",
46273=>X"00",
46274=>X"00",
46275=>X"00",
46276=>X"00",
46277=>X"00",
46278=>X"00",
46279=>X"00",
46280=>X"00",
46281=>X"00",
46282=>X"00",
46283=>X"00",
46284=>X"00",
46285=>X"00",
46286=>X"00",
46287=>X"00",
46288=>X"00",
46289=>X"00",
46290=>X"00",
46291=>X"00",
46292=>X"00",
46293=>X"00",
46294=>X"00",
46295=>X"00",
46296=>X"00",
46297=>X"00",
46298=>X"00",
46299=>X"00",
46300=>X"00",
46301=>X"00",
46302=>X"00",
46303=>X"00",
46304=>X"00",
46305=>X"00",
46306=>X"00",
46307=>X"00",
46308=>X"00",
46309=>X"00",
46310=>X"00",
46311=>X"00",
46312=>X"00",
46313=>X"00",
46314=>X"00",
46315=>X"00",
46316=>X"00",
46317=>X"00",
46318=>X"00",
46319=>X"00",
46320=>X"00",
46321=>X"00",
46322=>X"00",
46323=>X"00",
46324=>X"00",
46325=>X"00",
46326=>X"00",
46327=>X"00",
46328=>X"00",
46329=>X"00",
46330=>X"00",
46331=>X"00",
46332=>X"00",
46333=>X"00",
46334=>X"00",
46335=>X"00",
46336=>X"00",
46337=>X"00",
46338=>X"00",
46339=>X"00",
46340=>X"00",
46341=>X"00",
46342=>X"00",
46343=>X"00",
46344=>X"00",
46345=>X"00",
46346=>X"00",
46347=>X"00",
46348=>X"00",
46349=>X"00",
46350=>X"00",
46351=>X"00",
46352=>X"00",
46353=>X"00",
46354=>X"00",
46355=>X"00",
46356=>X"00",
46357=>X"00",
46358=>X"00",
46359=>X"00",
46360=>X"00",
46361=>X"00",
46362=>X"00",
46363=>X"00",
46364=>X"00",
46365=>X"00",
46366=>X"00",
46367=>X"00",
46368=>X"00",
46369=>X"00",
46370=>X"00",
46371=>X"00",
46372=>X"00",
46373=>X"00",
46374=>X"00",
46375=>X"00",
46376=>X"00",
46377=>X"00",
46378=>X"00",
46379=>X"00",
46380=>X"00",
46381=>X"00",
46382=>X"00",
46383=>X"00",
46384=>X"00",
46385=>X"00",
46386=>X"00",
46387=>X"00",
46388=>X"00",
46389=>X"00",
46390=>X"00",
46391=>X"00",
46392=>X"00",
46393=>X"00",
46394=>X"00",
46395=>X"00",
46396=>X"00",
46397=>X"00",
46398=>X"00",
46399=>X"00",
46400=>X"00",
46401=>X"00",
46402=>X"00",
46403=>X"00",
46404=>X"00",
46405=>X"00",
46406=>X"00",
46407=>X"00",
46408=>X"00",
46409=>X"00",
46410=>X"00",
46411=>X"00",
46412=>X"00",
46413=>X"00",
46414=>X"00",
46415=>X"00",
46416=>X"00",
46417=>X"00",
46418=>X"00",
46419=>X"00",
46420=>X"00",
46421=>X"00",
46422=>X"00",
46423=>X"00",
46424=>X"00",
46425=>X"00",
46426=>X"00",
46427=>X"00",
46428=>X"00",
46429=>X"00",
46430=>X"00",
46431=>X"00",
46432=>X"00",
46433=>X"00",
46434=>X"00",
46435=>X"00",
46436=>X"00",
46437=>X"00",
46438=>X"00",
46439=>X"00",
46440=>X"00",
46441=>X"00",
46442=>X"00",
46443=>X"00",
46444=>X"00",
46445=>X"00",
46446=>X"00",
46447=>X"00",
46448=>X"00",
46449=>X"00",
46450=>X"00",
46451=>X"00",
46452=>X"00",
46453=>X"00",
46454=>X"00",
46455=>X"00",
46456=>X"00",
46457=>X"00",
46458=>X"00",
46459=>X"00",
46460=>X"00",
46461=>X"00",
46462=>X"00",
46463=>X"00",
46464=>X"00",
46465=>X"00",
46466=>X"00",
46467=>X"00",
46468=>X"00",
46469=>X"00",
46470=>X"00",
46471=>X"00",
46472=>X"00",
46473=>X"00",
46474=>X"00",
46475=>X"00",
46476=>X"00",
46477=>X"00",
46478=>X"00",
46479=>X"00",
46480=>X"00",
46481=>X"00",
46482=>X"00",
46483=>X"00",
46484=>X"00",
46485=>X"00",
46486=>X"00",
46487=>X"00",
46488=>X"00",
46489=>X"00",
46490=>X"00",
46491=>X"00",
46492=>X"00",
46493=>X"00",
46494=>X"00",
46495=>X"00",
46496=>X"00",
46497=>X"00",
46498=>X"00",
46499=>X"00",
46500=>X"00",
46501=>X"00",
46502=>X"00",
46503=>X"00",
46504=>X"00",
46505=>X"00",
46506=>X"00",
46507=>X"00",
46508=>X"00",
46509=>X"00",
46510=>X"00",
46511=>X"00",
46512=>X"00",
46513=>X"00",
46514=>X"00",
46515=>X"00",
46516=>X"00",
46517=>X"00",
46518=>X"00",
46519=>X"00",
46520=>X"00",
46521=>X"00",
46522=>X"00",
46523=>X"00",
46524=>X"00",
46525=>X"00",
46526=>X"00",
46527=>X"00",
46528=>X"00",
46529=>X"00",
46530=>X"00",
46531=>X"00",
46532=>X"00",
46533=>X"00",
46534=>X"00",
46535=>X"00",
46536=>X"00",
46537=>X"00",
46538=>X"00",
46539=>X"00",
46540=>X"00",
46541=>X"00",
46542=>X"00",
46543=>X"00",
46544=>X"00",
46545=>X"00",
46546=>X"00",
46547=>X"00",
46548=>X"00",
46549=>X"00",
46550=>X"00",
46551=>X"00",
46552=>X"00",
46553=>X"00",
46554=>X"00",
46555=>X"00",
46556=>X"00",
46557=>X"00",
46558=>X"00",
46559=>X"00",
46560=>X"00",
46561=>X"00",
46562=>X"00",
46563=>X"00",
46564=>X"00",
46565=>X"00",
46566=>X"00",
46567=>X"00",
46568=>X"00",
46569=>X"00",
46570=>X"00",
46571=>X"00",
46572=>X"00",
46573=>X"00",
46574=>X"00",
46575=>X"00",
46576=>X"00",
46577=>X"00",
46578=>X"00",
46579=>X"00",
46580=>X"00",
46581=>X"00",
46582=>X"00",
46583=>X"00",
46584=>X"00",
46585=>X"00",
46586=>X"00",
46587=>X"00",
46588=>X"00",
46589=>X"00",
46590=>X"00",
46591=>X"00",
46592=>X"00",
46593=>X"00",
46594=>X"00",
46595=>X"00",
46596=>X"00",
46597=>X"00",
46598=>X"00",
46599=>X"00",
46600=>X"00",
46601=>X"00",
46602=>X"00",
46603=>X"00",
46604=>X"00",
46605=>X"00",
46606=>X"00",
46607=>X"00",
46608=>X"00",
46609=>X"00",
46610=>X"00",
46611=>X"00",
46612=>X"00",
46613=>X"00",
46614=>X"00",
46615=>X"00",
46616=>X"00",
46617=>X"00",
46618=>X"00",
46619=>X"00",
46620=>X"00",
46621=>X"00",
46622=>X"00",
46623=>X"00",
46624=>X"00",
46625=>X"00",
46626=>X"00",
46627=>X"00",
46628=>X"00",
46629=>X"00",
46630=>X"00",
46631=>X"00",
46632=>X"00",
46633=>X"00",
46634=>X"00",
46635=>X"00",
46636=>X"00",
46637=>X"00",
46638=>X"00",
46639=>X"00",
46640=>X"00",
46641=>X"00",
46642=>X"00",
46643=>X"00",
46644=>X"00",
46645=>X"00",
46646=>X"00",
46647=>X"00",
46648=>X"00",
46649=>X"00",
46650=>X"00",
46651=>X"00",
46652=>X"00",
46653=>X"00",
46654=>X"00",
46655=>X"00",
46656=>X"00",
46657=>X"00",
46658=>X"00",
46659=>X"00",
46660=>X"00",
46661=>X"00",
46662=>X"00",
46663=>X"00",
46664=>X"00",
46665=>X"00",
46666=>X"00",
46667=>X"00",
46668=>X"00",
46669=>X"00",
46670=>X"00",
46671=>X"00",
46672=>X"00",
46673=>X"00",
46674=>X"00",
46675=>X"00",
46676=>X"00",
46677=>X"00",
46678=>X"00",
46679=>X"00",
46680=>X"00",
46681=>X"00",
46682=>X"00",
46683=>X"00",
46684=>X"00",
46685=>X"00",
46686=>X"00",
46687=>X"00",
46688=>X"00",
46689=>X"00",
46690=>X"00",
46691=>X"00",
46692=>X"00",
46693=>X"00",
46694=>X"00",
46695=>X"00",
46696=>X"00",
46697=>X"00",
46698=>X"00",
46699=>X"00",
46700=>X"00",
46701=>X"00",
46702=>X"00",
46703=>X"00",
46704=>X"00",
46705=>X"00",
46706=>X"00",
46707=>X"00",
46708=>X"00",
46709=>X"00",
46710=>X"00",
46711=>X"00",
46712=>X"00",
46713=>X"00",
46714=>X"00",
46715=>X"00",
46716=>X"00",
46717=>X"00",
46718=>X"00",
46719=>X"00",
46720=>X"00",
46721=>X"00",
46722=>X"00",
46723=>X"00",
46724=>X"00",
46725=>X"00",
46726=>X"00",
46727=>X"00",
46728=>X"00",
46729=>X"00",
46730=>X"00",
46731=>X"00",
46732=>X"00",
46733=>X"00",
46734=>X"00",
46735=>X"00",
46736=>X"00",
46737=>X"00",
46738=>X"00",
46739=>X"00",
46740=>X"00",
46741=>X"00",
46742=>X"00",
46743=>X"00",
46744=>X"00",
46745=>X"00",
46746=>X"00",
46747=>X"00",
46748=>X"00",
46749=>X"00",
46750=>X"00",
46751=>X"00",
46752=>X"00",
46753=>X"00",
46754=>X"00",
46755=>X"00",
46756=>X"00",
46757=>X"00",
46758=>X"00",
46759=>X"00",
46760=>X"00",
46761=>X"00",
46762=>X"00",
46763=>X"00",
46764=>X"00",
46765=>X"00",
46766=>X"00",
46767=>X"00",
46768=>X"00",
46769=>X"00",
46770=>X"00",
46771=>X"00",
46772=>X"00",
46773=>X"00",
46774=>X"00",
46775=>X"00",
46776=>X"00",
46777=>X"00",
46778=>X"00",
46779=>X"00",
46780=>X"00",
46781=>X"00",
46782=>X"00",
46783=>X"00",
46784=>X"00",
46785=>X"00",
46786=>X"00",
46787=>X"00",
46788=>X"00",
46789=>X"00",
46790=>X"00",
46791=>X"00",
46792=>X"00",
46793=>X"00",
46794=>X"00",
46795=>X"00",
46796=>X"00",
46797=>X"00",
46798=>X"00",
46799=>X"00",
46800=>X"00",
46801=>X"00",
46802=>X"00",
46803=>X"00",
46804=>X"00",
46805=>X"00",
46806=>X"00",
46807=>X"00",
46808=>X"00",
46809=>X"00",
46810=>X"00",
46811=>X"00",
46812=>X"00",
46813=>X"00",
46814=>X"00",
46815=>X"00",
46816=>X"00",
46817=>X"00",
46818=>X"00",
46819=>X"00",
46820=>X"00",
46821=>X"00",
46822=>X"00",
46823=>X"00",
46824=>X"00",
46825=>X"00",
46826=>X"00",
46827=>X"00",
46828=>X"00",
46829=>X"00",
46830=>X"00",
46831=>X"00",
46832=>X"00",
46833=>X"00",
46834=>X"00",
46835=>X"00",
46836=>X"00",
46837=>X"00",
46838=>X"00",
46839=>X"00",
46840=>X"00",
46841=>X"00",
46842=>X"00",
46843=>X"00",
46844=>X"00",
46845=>X"00",
46846=>X"00",
46847=>X"00",
46848=>X"00",
46849=>X"00",
46850=>X"00",
46851=>X"00",
46852=>X"00",
46853=>X"00",
46854=>X"00",
46855=>X"00",
46856=>X"00",
46857=>X"00",
46858=>X"00",
46859=>X"00",
46860=>X"00",
46861=>X"00",
46862=>X"00",
46863=>X"00",
46864=>X"00",
46865=>X"00",
46866=>X"00",
46867=>X"00",
46868=>X"00",
46869=>X"00",
46870=>X"00",
46871=>X"00",
46872=>X"00",
46873=>X"00",
46874=>X"00",
46875=>X"00",
46876=>X"00",
46877=>X"00",
46878=>X"00",
46879=>X"00",
46880=>X"00",
46881=>X"00",
46882=>X"00",
46883=>X"00",
46884=>X"00",
46885=>X"00",
46886=>X"00",
46887=>X"00",
46888=>X"00",
46889=>X"00",
46890=>X"00",
46891=>X"00",
46892=>X"00",
46893=>X"00",
46894=>X"00",
46895=>X"00",
46896=>X"00",
46897=>X"00",
46898=>X"00",
46899=>X"00",
46900=>X"00",
46901=>X"00",
46902=>X"00",
46903=>X"00",
46904=>X"00",
46905=>X"00",
46906=>X"00",
46907=>X"00",
46908=>X"00",
46909=>X"00",
46910=>X"00",
46911=>X"00",
46912=>X"00",
46913=>X"00",
46914=>X"00",
46915=>X"00",
46916=>X"00",
46917=>X"00",
46918=>X"00",
46919=>X"00",
46920=>X"00",
46921=>X"00",
46922=>X"00",
46923=>X"00",
46924=>X"00",
46925=>X"00",
46926=>X"00",
46927=>X"00",
46928=>X"00",
46929=>X"00",
46930=>X"00",
46931=>X"00",
46932=>X"00",
46933=>X"00",
46934=>X"00",
46935=>X"00",
46936=>X"00",
46937=>X"00",
46938=>X"00",
46939=>X"00",
46940=>X"00",
46941=>X"00",
46942=>X"00",
46943=>X"00",
46944=>X"00",
46945=>X"00",
46946=>X"00",
46947=>X"00",
46948=>X"00",
46949=>X"00",
46950=>X"00",
46951=>X"00",
46952=>X"00",
46953=>X"00",
46954=>X"00",
46955=>X"00",
46956=>X"00",
46957=>X"00",
46958=>X"00",
46959=>X"00",
46960=>X"00",
46961=>X"00",
46962=>X"00",
46963=>X"00",
46964=>X"00",
46965=>X"00",
46966=>X"00",
46967=>X"00",
46968=>X"00",
46969=>X"00",
46970=>X"00",
46971=>X"00",
46972=>X"00",
46973=>X"00",
46974=>X"00",
46975=>X"00",
46976=>X"00",
46977=>X"00",
46978=>X"00",
46979=>X"00",
46980=>X"00",
46981=>X"00",
46982=>X"00",
46983=>X"00",
46984=>X"00",
46985=>X"00",
46986=>X"00",
46987=>X"00",
46988=>X"00",
46989=>X"00",
46990=>X"00",
46991=>X"00",
46992=>X"00",
46993=>X"00",
46994=>X"00",
46995=>X"00",
46996=>X"00",
46997=>X"00",
46998=>X"00",
46999=>X"00",
47000=>X"00",
47001=>X"00",
47002=>X"00",
47003=>X"00",
47004=>X"00",
47005=>X"00",
47006=>X"00",
47007=>X"00",
47008=>X"00",
47009=>X"00",
47010=>X"00",
47011=>X"00",
47012=>X"00",
47013=>X"00",
47014=>X"00",
47015=>X"00",
47016=>X"00",
47017=>X"00",
47018=>X"00",
47019=>X"00",
47020=>X"00",
47021=>X"00",
47022=>X"00",
47023=>X"00",
47024=>X"00",
47025=>X"00",
47026=>X"00",
47027=>X"00",
47028=>X"00",
47029=>X"00",
47030=>X"00",
47031=>X"00",
47032=>X"00",
47033=>X"00",
47034=>X"00",
47035=>X"00",
47036=>X"00",
47037=>X"00",
47038=>X"00",
47039=>X"00",
47040=>X"00",
47041=>X"00",
47042=>X"00",
47043=>X"00",
47044=>X"00",
47045=>X"00",
47046=>X"00",
47047=>X"00",
47048=>X"00",
47049=>X"00",
47050=>X"00",
47051=>X"00",
47052=>X"00",
47053=>X"00",
47054=>X"00",
47055=>X"00",
47056=>X"00",
47057=>X"00",
47058=>X"00",
47059=>X"00",
47060=>X"00",
47061=>X"00",
47062=>X"00",
47063=>X"00",
47064=>X"00",
47065=>X"00",
47066=>X"00",
47067=>X"00",
47068=>X"00",
47069=>X"00",
47070=>X"00",
47071=>X"00",
47072=>X"00",
47073=>X"00",
47074=>X"00",
47075=>X"00",
47076=>X"00",
47077=>X"00",
47078=>X"00",
47079=>X"00",
47080=>X"00",
47081=>X"00",
47082=>X"00",
47083=>X"00",
47084=>X"00",
47085=>X"00",
47086=>X"00",
47087=>X"00",
47088=>X"00",
47089=>X"00",
47090=>X"00",
47091=>X"00",
47092=>X"00",
47093=>X"00",
47094=>X"00",
47095=>X"00",
47096=>X"00",
47097=>X"00",
47098=>X"00",
47099=>X"00",
47100=>X"00",
47101=>X"00",
47102=>X"00",
47103=>X"00",
47104=>X"00",
47105=>X"00",
47106=>X"00",
47107=>X"00",
47108=>X"00",
47109=>X"00",
47110=>X"00",
47111=>X"00",
47112=>X"00",
47113=>X"00",
47114=>X"00",
47115=>X"00",
47116=>X"00",
47117=>X"00",
47118=>X"00",
47119=>X"00",
47120=>X"00",
47121=>X"00",
47122=>X"00",
47123=>X"00",
47124=>X"00",
47125=>X"00",
47126=>X"00",
47127=>X"00",
47128=>X"00",
47129=>X"00",
47130=>X"00",
47131=>X"00",
47132=>X"00",
47133=>X"00",
47134=>X"00",
47135=>X"00",
47136=>X"00",
47137=>X"00",
47138=>X"00",
47139=>X"00",
47140=>X"00",
47141=>X"00",
47142=>X"00",
47143=>X"00",
47144=>X"00",
47145=>X"00",
47146=>X"00",
47147=>X"00",
47148=>X"00",
47149=>X"00",
47150=>X"00",
47151=>X"00",
47152=>X"00",
47153=>X"00",
47154=>X"00",
47155=>X"00",
47156=>X"00",
47157=>X"00",
47158=>X"00",
47159=>X"00",
47160=>X"00",
47161=>X"00",
47162=>X"00",
47163=>X"00",
47164=>X"00",
47165=>X"00",
47166=>X"00",
47167=>X"00",
47168=>X"00",
47169=>X"00",
47170=>X"00",
47171=>X"00",
47172=>X"00",
47173=>X"00",
47174=>X"00",
47175=>X"00",
47176=>X"00",
47177=>X"00",
47178=>X"00",
47179=>X"00",
47180=>X"00",
47181=>X"00",
47182=>X"00",
47183=>X"00",
47184=>X"00",
47185=>X"00",
47186=>X"00",
47187=>X"00",
47188=>X"00",
47189=>X"00",
47190=>X"00",
47191=>X"00",
47192=>X"00",
47193=>X"00",
47194=>X"00",
47195=>X"00",
47196=>X"00",
47197=>X"00",
47198=>X"00",
47199=>X"00",
47200=>X"00",
47201=>X"00",
47202=>X"00",
47203=>X"00",
47204=>X"00",
47205=>X"00",
47206=>X"00",
47207=>X"00",
47208=>X"00",
47209=>X"00",
47210=>X"00",
47211=>X"00",
47212=>X"00",
47213=>X"00",
47214=>X"00",
47215=>X"00",
47216=>X"00",
47217=>X"00",
47218=>X"00",
47219=>X"00",
47220=>X"00",
47221=>X"00",
47222=>X"00",
47223=>X"00",
47224=>X"00",
47225=>X"00",
47226=>X"00",
47227=>X"00",
47228=>X"00",
47229=>X"00",
47230=>X"00",
47231=>X"00",
47232=>X"00",
47233=>X"00",
47234=>X"00",
47235=>X"00",
47236=>X"00",
47237=>X"00",
47238=>X"00",
47239=>X"00",
47240=>X"00",
47241=>X"00",
47242=>X"00",
47243=>X"00",
47244=>X"00",
47245=>X"00",
47246=>X"00",
47247=>X"00",
47248=>X"00",
47249=>X"00",
47250=>X"00",
47251=>X"00",
47252=>X"00",
47253=>X"00",
47254=>X"00",
47255=>X"00",
47256=>X"00",
47257=>X"00",
47258=>X"00",
47259=>X"00",
47260=>X"00",
47261=>X"00",
47262=>X"00",
47263=>X"00",
47264=>X"00",
47265=>X"00",
47266=>X"00",
47267=>X"00",
47268=>X"00",
47269=>X"00",
47270=>X"00",
47271=>X"00",
47272=>X"00",
47273=>X"00",
47274=>X"00",
47275=>X"00",
47276=>X"00",
47277=>X"00",
47278=>X"00",
47279=>X"00",
47280=>X"00",
47281=>X"00",
47282=>X"00",
47283=>X"00",
47284=>X"00",
47285=>X"00",
47286=>X"00",
47287=>X"00",
47288=>X"00",
47289=>X"00",
47290=>X"00",
47291=>X"00",
47292=>X"00",
47293=>X"00",
47294=>X"00",
47295=>X"00",
47296=>X"00",
47297=>X"00",
47298=>X"00",
47299=>X"00",
47300=>X"00",
47301=>X"00",
47302=>X"00",
47303=>X"00",
47304=>X"00",
47305=>X"00",
47306=>X"00",
47307=>X"00",
47308=>X"00",
47309=>X"00",
47310=>X"00",
47311=>X"00",
47312=>X"00",
47313=>X"00",
47314=>X"00",
47315=>X"00",
47316=>X"00",
47317=>X"00",
47318=>X"00",
47319=>X"00",
47320=>X"00",
47321=>X"00",
47322=>X"00",
47323=>X"00",
47324=>X"00",
47325=>X"00",
47326=>X"00",
47327=>X"00",
47328=>X"00",
47329=>X"00",
47330=>X"00",
47331=>X"00",
47332=>X"00",
47333=>X"00",
47334=>X"00",
47335=>X"00",
47336=>X"00",
47337=>X"00",
47338=>X"00",
47339=>X"00",
47340=>X"00",
47341=>X"00",
47342=>X"00",
47343=>X"00",
47344=>X"00",
47345=>X"00",
47346=>X"00",
47347=>X"00",
47348=>X"00",
47349=>X"00",
47350=>X"00",
47351=>X"00",
47352=>X"00",
47353=>X"00",
47354=>X"00",
47355=>X"00",
47356=>X"00",
47357=>X"00",
47358=>X"00",
47359=>X"00",
47360=>X"00",
47361=>X"00",
47362=>X"00",
47363=>X"00",
47364=>X"00",
47365=>X"00",
47366=>X"00",
47367=>X"00",
47368=>X"00",
47369=>X"00",
47370=>X"00",
47371=>X"00",
47372=>X"00",
47373=>X"00",
47374=>X"00",
47375=>X"00",
47376=>X"00",
47377=>X"00",
47378=>X"00",
47379=>X"00",
47380=>X"00",
47381=>X"00",
47382=>X"00",
47383=>X"00",
47384=>X"00",
47385=>X"00",
47386=>X"00",
47387=>X"00",
47388=>X"00",
47389=>X"00",
47390=>X"00",
47391=>X"00",
47392=>X"00",
47393=>X"00",
47394=>X"00",
47395=>X"00",
47396=>X"00",
47397=>X"00",
47398=>X"00",
47399=>X"00",
47400=>X"00",
47401=>X"00",
47402=>X"00",
47403=>X"00",
47404=>X"00",
47405=>X"00",
47406=>X"00",
47407=>X"00",
47408=>X"00",
47409=>X"00",
47410=>X"00",
47411=>X"00",
47412=>X"00",
47413=>X"00",
47414=>X"00",
47415=>X"00",
47416=>X"00",
47417=>X"00",
47418=>X"00",
47419=>X"00",
47420=>X"00",
47421=>X"00",
47422=>X"00",
47423=>X"00",
47424=>X"00",
47425=>X"00",
47426=>X"00",
47427=>X"00",
47428=>X"00",
47429=>X"00",
47430=>X"00",
47431=>X"00",
47432=>X"00",
47433=>X"00",
47434=>X"00",
47435=>X"00",
47436=>X"00",
47437=>X"00",
47438=>X"00",
47439=>X"00",
47440=>X"00",
47441=>X"00",
47442=>X"00",
47443=>X"00",
47444=>X"00",
47445=>X"00",
47446=>X"00",
47447=>X"00",
47448=>X"00",
47449=>X"00",
47450=>X"00",
47451=>X"00",
47452=>X"00",
47453=>X"00",
47454=>X"00",
47455=>X"00",
47456=>X"00",
47457=>X"00",
47458=>X"00",
47459=>X"00",
47460=>X"00",
47461=>X"00",
47462=>X"00",
47463=>X"00",
47464=>X"00",
47465=>X"00",
47466=>X"00",
47467=>X"00",
47468=>X"00",
47469=>X"00",
47470=>X"00",
47471=>X"00",
47472=>X"00",
47473=>X"00",
47474=>X"00",
47475=>X"00",
47476=>X"00",
47477=>X"00",
47478=>X"00",
47479=>X"00",
47480=>X"00",
47481=>X"00",
47482=>X"00",
47483=>X"00",
47484=>X"00",
47485=>X"00",
47486=>X"00",
47487=>X"00",
47488=>X"00",
47489=>X"00",
47490=>X"00",
47491=>X"00",
47492=>X"00",
47493=>X"00",
47494=>X"00",
47495=>X"00",
47496=>X"00",
47497=>X"00",
47498=>X"00",
47499=>X"00",
47500=>X"00",
47501=>X"00",
47502=>X"00",
47503=>X"00",
47504=>X"00",
47505=>X"00",
47506=>X"00",
47507=>X"00",
47508=>X"00",
47509=>X"00",
47510=>X"00",
47511=>X"00",
47512=>X"00",
47513=>X"00",
47514=>X"00",
47515=>X"00",
47516=>X"00",
47517=>X"00",
47518=>X"00",
47519=>X"00",
47520=>X"00",
47521=>X"00",
47522=>X"00",
47523=>X"00",
47524=>X"00",
47525=>X"00",
47526=>X"00",
47527=>X"00",
47528=>X"00",
47529=>X"00",
47530=>X"00",
47531=>X"00",
47532=>X"00",
47533=>X"00",
47534=>X"00",
47535=>X"00",
47536=>X"00",
47537=>X"00",
47538=>X"00",
47539=>X"00",
47540=>X"00",
47541=>X"00",
47542=>X"00",
47543=>X"00",
47544=>X"00",
47545=>X"00",
47546=>X"00",
47547=>X"00",
47548=>X"00",
47549=>X"00",
47550=>X"00",
47551=>X"00",
47552=>X"00",
47553=>X"00",
47554=>X"00",
47555=>X"00",
47556=>X"00",
47557=>X"00",
47558=>X"00",
47559=>X"00",
47560=>X"00",
47561=>X"00",
47562=>X"00",
47563=>X"00",
47564=>X"00",
47565=>X"00",
47566=>X"00",
47567=>X"00",
47568=>X"00",
47569=>X"00",
47570=>X"00",
47571=>X"00",
47572=>X"00",
47573=>X"00",
47574=>X"00",
47575=>X"00",
47576=>X"00",
47577=>X"00",
47578=>X"00",
47579=>X"00",
47580=>X"00",
47581=>X"00",
47582=>X"00",
47583=>X"00",
47584=>X"00",
47585=>X"00",
47586=>X"00",
47587=>X"00",
47588=>X"00",
47589=>X"00",
47590=>X"00",
47591=>X"00",
47592=>X"00",
47593=>X"00",
47594=>X"00",
47595=>X"00",
47596=>X"00",
47597=>X"00",
47598=>X"00",
47599=>X"00",
47600=>X"00",
47601=>X"00",
47602=>X"00",
47603=>X"00",
47604=>X"00",
47605=>X"00",
47606=>X"00",
47607=>X"00",
47608=>X"00",
47609=>X"00",
47610=>X"00",
47611=>X"00",
47612=>X"00",
47613=>X"00",
47614=>X"00",
47615=>X"00",
47616=>X"00",
47617=>X"00",
47618=>X"00",
47619=>X"00",
47620=>X"00",
47621=>X"00",
47622=>X"00",
47623=>X"00",
47624=>X"00",
47625=>X"00",
47626=>X"00",
47627=>X"00",
47628=>X"00",
47629=>X"00",
47630=>X"00",
47631=>X"00",
47632=>X"00",
47633=>X"00",
47634=>X"00",
47635=>X"00",
47636=>X"00",
47637=>X"00",
47638=>X"00",
47639=>X"00",
47640=>X"00",
47641=>X"00",
47642=>X"00",
47643=>X"00",
47644=>X"00",
47645=>X"00",
47646=>X"00",
47647=>X"00",
47648=>X"00",
47649=>X"00",
47650=>X"00",
47651=>X"00",
47652=>X"00",
47653=>X"00",
47654=>X"00",
47655=>X"00",
47656=>X"00",
47657=>X"00",
47658=>X"00",
47659=>X"00",
47660=>X"00",
47661=>X"00",
47662=>X"00",
47663=>X"00",
47664=>X"00",
47665=>X"00",
47666=>X"00",
47667=>X"00",
47668=>X"00",
47669=>X"00",
47670=>X"00",
47671=>X"00",
47672=>X"00",
47673=>X"00",
47674=>X"00",
47675=>X"00",
47676=>X"00",
47677=>X"00",
47678=>X"00",
47679=>X"00",
47680=>X"00",
47681=>X"00",
47682=>X"00",
47683=>X"00",
47684=>X"00",
47685=>X"00",
47686=>X"00",
47687=>X"00",
47688=>X"00",
47689=>X"00",
47690=>X"00",
47691=>X"00",
47692=>X"00",
47693=>X"00",
47694=>X"00",
47695=>X"00",
47696=>X"00",
47697=>X"00",
47698=>X"00",
47699=>X"00",
47700=>X"00",
47701=>X"00",
47702=>X"00",
47703=>X"00",
47704=>X"00",
47705=>X"00",
47706=>X"00",
47707=>X"00",
47708=>X"00",
47709=>X"00",
47710=>X"00",
47711=>X"00",
47712=>X"00",
47713=>X"00",
47714=>X"00",
47715=>X"00",
47716=>X"00",
47717=>X"00",
47718=>X"00",
47719=>X"00",
47720=>X"00",
47721=>X"00",
47722=>X"00",
47723=>X"00",
47724=>X"00",
47725=>X"00",
47726=>X"00",
47727=>X"00",
47728=>X"00",
47729=>X"00",
47730=>X"00",
47731=>X"00",
47732=>X"00",
47733=>X"00",
47734=>X"00",
47735=>X"00",
47736=>X"00",
47737=>X"00",
47738=>X"00",
47739=>X"00",
47740=>X"00",
47741=>X"00",
47742=>X"00",
47743=>X"00",
47744=>X"00",
47745=>X"00",
47746=>X"00",
47747=>X"00",
47748=>X"00",
47749=>X"00",
47750=>X"00",
47751=>X"00",
47752=>X"00",
47753=>X"00",
47754=>X"00",
47755=>X"00",
47756=>X"00",
47757=>X"00",
47758=>X"00",
47759=>X"00",
47760=>X"00",
47761=>X"00",
47762=>X"00",
47763=>X"00",
47764=>X"00",
47765=>X"00",
47766=>X"00",
47767=>X"00",
47768=>X"00",
47769=>X"00",
47770=>X"00",
47771=>X"00",
47772=>X"00",
47773=>X"00",
47774=>X"00",
47775=>X"00",
47776=>X"00",
47777=>X"00",
47778=>X"00",
47779=>X"00",
47780=>X"00",
47781=>X"00",
47782=>X"00",
47783=>X"00",
47784=>X"00",
47785=>X"00",
47786=>X"00",
47787=>X"00",
47788=>X"00",
47789=>X"00",
47790=>X"00",
47791=>X"00",
47792=>X"00",
47793=>X"00",
47794=>X"00",
47795=>X"00",
47796=>X"00",
47797=>X"00",
47798=>X"00",
47799=>X"00",
47800=>X"00",
47801=>X"00",
47802=>X"00",
47803=>X"00",
47804=>X"00",
47805=>X"00",
47806=>X"00",
47807=>X"00",
47808=>X"00",
47809=>X"00",
47810=>X"00",
47811=>X"00",
47812=>X"00",
47813=>X"00",
47814=>X"00",
47815=>X"00",
47816=>X"00",
47817=>X"00",
47818=>X"00",
47819=>X"00",
47820=>X"00",
47821=>X"00",
47822=>X"00",
47823=>X"00",
47824=>X"00",
47825=>X"00",
47826=>X"00",
47827=>X"00",
47828=>X"00",
47829=>X"00",
47830=>X"00",
47831=>X"00",
47832=>X"00",
47833=>X"00",
47834=>X"00",
47835=>X"00",
47836=>X"00",
47837=>X"00",
47838=>X"00",
47839=>X"00",
47840=>X"00",
47841=>X"00",
47842=>X"00",
47843=>X"00",
47844=>X"00",
47845=>X"00",
47846=>X"00",
47847=>X"00",
47848=>X"00",
47849=>X"00",
47850=>X"00",
47851=>X"00",
47852=>X"00",
47853=>X"00",
47854=>X"00",
47855=>X"00",
47856=>X"00",
47857=>X"00",
47858=>X"00",
47859=>X"00",
47860=>X"00",
47861=>X"00",
47862=>X"00",
47863=>X"00",
47864=>X"00",
47865=>X"00",
47866=>X"00",
47867=>X"00",
47868=>X"00",
47869=>X"00",
47870=>X"00",
47871=>X"00",
47872=>X"00",
47873=>X"00",
47874=>X"00",
47875=>X"00",
47876=>X"00",
47877=>X"00",
47878=>X"00",
47879=>X"00",
47880=>X"00",
47881=>X"00",
47882=>X"00",
47883=>X"00",
47884=>X"00",
47885=>X"00",
47886=>X"00",
47887=>X"00",
47888=>X"00",
47889=>X"00",
47890=>X"00",
47891=>X"00",
47892=>X"00",
47893=>X"00",
47894=>X"00",
47895=>X"00",
47896=>X"00",
47897=>X"00",
47898=>X"00",
47899=>X"00",
47900=>X"00",
47901=>X"00",
47902=>X"00",
47903=>X"00",
47904=>X"00",
47905=>X"00",
47906=>X"00",
47907=>X"00",
47908=>X"00",
47909=>X"00",
47910=>X"00",
47911=>X"00",
47912=>X"00",
47913=>X"00",
47914=>X"00",
47915=>X"00",
47916=>X"00",
47917=>X"00",
47918=>X"00",
47919=>X"00",
47920=>X"00",
47921=>X"00",
47922=>X"00",
47923=>X"00",
47924=>X"00",
47925=>X"00",
47926=>X"00",
47927=>X"00",
47928=>X"00",
47929=>X"00",
47930=>X"00",
47931=>X"00",
47932=>X"00",
47933=>X"00",
47934=>X"00",
47935=>X"00",
47936=>X"00",
47937=>X"00",
47938=>X"00",
47939=>X"00",
47940=>X"00",
47941=>X"00",
47942=>X"00",
47943=>X"00",
47944=>X"00",
47945=>X"00",
47946=>X"00",
47947=>X"00",
47948=>X"00",
47949=>X"00",
47950=>X"00",
47951=>X"00",
47952=>X"00",
47953=>X"00",
47954=>X"00",
47955=>X"00",
47956=>X"00",
47957=>X"00",
47958=>X"00",
47959=>X"00",
47960=>X"00",
47961=>X"00",
47962=>X"00",
47963=>X"00",
47964=>X"00",
47965=>X"00",
47966=>X"00",
47967=>X"00",
47968=>X"00",
47969=>X"00",
47970=>X"00",
47971=>X"00",
47972=>X"00",
47973=>X"00",
47974=>X"00",
47975=>X"00",
47976=>X"00",
47977=>X"00",
47978=>X"00",
47979=>X"00",
47980=>X"00",
47981=>X"00",
47982=>X"00",
47983=>X"00",
47984=>X"00",
47985=>X"00",
47986=>X"00",
47987=>X"00",
47988=>X"00",
47989=>X"00",
47990=>X"00",
47991=>X"00",
47992=>X"00",
47993=>X"00",
47994=>X"00",
47995=>X"00",
47996=>X"00",
47997=>X"00",
47998=>X"00",
47999=>X"00",
48000=>X"00",
48001=>X"00",
48002=>X"00",
48003=>X"00",
48004=>X"00",
48005=>X"00",
48006=>X"00",
48007=>X"00",
48008=>X"00",
48009=>X"00",
48010=>X"00",
48011=>X"00",
48012=>X"00",
48013=>X"00",
48014=>X"00",
48015=>X"00",
48016=>X"00",
48017=>X"00",
48018=>X"00",
48019=>X"00",
48020=>X"00",
48021=>X"00",
48022=>X"00",
48023=>X"00",
48024=>X"00",
48025=>X"00",
48026=>X"00",
48027=>X"00",
48028=>X"00",
48029=>X"00",
48030=>X"00",
48031=>X"00",
48032=>X"00",
48033=>X"00",
48034=>X"00",
48035=>X"00",
48036=>X"00",
48037=>X"00",
48038=>X"00",
48039=>X"00",
48040=>X"00",
48041=>X"00",
48042=>X"00",
48043=>X"00",
48044=>X"00",
48045=>X"00",
48046=>X"00",
48047=>X"00",
48048=>X"00",
48049=>X"00",
48050=>X"00",
48051=>X"00",
48052=>X"00",
48053=>X"00",
48054=>X"00",
48055=>X"00",
48056=>X"00",
48057=>X"00",
48058=>X"00",
48059=>X"00",
48060=>X"00",
48061=>X"00",
48062=>X"00",
48063=>X"00",
48064=>X"00",
48065=>X"00",
48066=>X"00",
48067=>X"00",
48068=>X"00",
48069=>X"00",
48070=>X"00",
48071=>X"00",
48072=>X"00",
48073=>X"00",
48074=>X"00",
48075=>X"00",
48076=>X"00",
48077=>X"00",
48078=>X"00",
48079=>X"00",
48080=>X"00",
48081=>X"00",
48082=>X"00",
48083=>X"00",
48084=>X"00",
48085=>X"00",
48086=>X"00",
48087=>X"00",
48088=>X"00",
48089=>X"00",
48090=>X"00",
48091=>X"00",
48092=>X"00",
48093=>X"00",
48094=>X"00",
48095=>X"00",
48096=>X"00",
48097=>X"00",
48098=>X"00",
48099=>X"00",
48100=>X"00",
48101=>X"00",
48102=>X"00",
48103=>X"00",
48104=>X"00",
48105=>X"00",
48106=>X"00",
48107=>X"00",
48108=>X"00",
48109=>X"00",
48110=>X"00",
48111=>X"00",
48112=>X"00",
48113=>X"00",
48114=>X"00",
48115=>X"00",
48116=>X"00",
48117=>X"00",
48118=>X"00",
48119=>X"00",
48120=>X"00",
48121=>X"00",
48122=>X"00",
48123=>X"00",
48124=>X"00",
48125=>X"00",
48126=>X"00",
48127=>X"00",
48128=>X"00",
48129=>X"00",
48130=>X"00",
48131=>X"00",
48132=>X"00",
48133=>X"00",
48134=>X"00",
48135=>X"00",
48136=>X"00",
48137=>X"00",
48138=>X"00",
48139=>X"00",
48140=>X"00",
48141=>X"00",
48142=>X"00",
48143=>X"00",
48144=>X"00",
48145=>X"00",
48146=>X"00",
48147=>X"00",
48148=>X"00",
48149=>X"00",
48150=>X"00",
48151=>X"00",
48152=>X"00",
48153=>X"00",
48154=>X"00",
48155=>X"00",
48156=>X"00",
48157=>X"00",
48158=>X"00",
48159=>X"00",
48160=>X"00",
48161=>X"00",
48162=>X"00",
48163=>X"00",
48164=>X"00",
48165=>X"00",
48166=>X"00",
48167=>X"00",
48168=>X"00",
48169=>X"00",
48170=>X"00",
48171=>X"00",
48172=>X"00",
48173=>X"00",
48174=>X"00",
48175=>X"00",
48176=>X"00",
48177=>X"00",
48178=>X"00",
48179=>X"00",
48180=>X"00",
48181=>X"00",
48182=>X"00",
48183=>X"00",
48184=>X"00",
48185=>X"00",
48186=>X"00",
48187=>X"00",
48188=>X"00",
48189=>X"00",
48190=>X"00",
48191=>X"00",
48192=>X"00",
48193=>X"00",
48194=>X"00",
48195=>X"00",
48196=>X"00",
48197=>X"00",
48198=>X"00",
48199=>X"00",
48200=>X"00",
48201=>X"00",
48202=>X"00",
48203=>X"00",
48204=>X"00",
48205=>X"00",
48206=>X"00",
48207=>X"00",
48208=>X"00",
48209=>X"00",
48210=>X"00",
48211=>X"00",
48212=>X"00",
48213=>X"00",
48214=>X"00",
48215=>X"00",
48216=>X"00",
48217=>X"00",
48218=>X"00",
48219=>X"00",
48220=>X"00",
48221=>X"00",
48222=>X"00",
48223=>X"00",
48224=>X"00",
48225=>X"00",
48226=>X"00",
48227=>X"00",
48228=>X"00",
48229=>X"00",
48230=>X"00",
48231=>X"00",
48232=>X"00",
48233=>X"00",
48234=>X"00",
48235=>X"00",
48236=>X"00",
48237=>X"00",
48238=>X"00",
48239=>X"00",
48240=>X"00",
48241=>X"00",
48242=>X"00",
48243=>X"00",
48244=>X"00",
48245=>X"00",
48246=>X"00",
48247=>X"00",
48248=>X"00",
48249=>X"00",
48250=>X"00",
48251=>X"00",
48252=>X"00",
48253=>X"00",
48254=>X"00",
48255=>X"00",
48256=>X"00",
48257=>X"00",
48258=>X"00",
48259=>X"00",
48260=>X"00",
48261=>X"00",
48262=>X"00",
48263=>X"00",
48264=>X"00",
48265=>X"00",
48266=>X"00",
48267=>X"00",
48268=>X"00",
48269=>X"00",
48270=>X"00",
48271=>X"00",
48272=>X"00",
48273=>X"00",
48274=>X"00",
48275=>X"00",
48276=>X"00",
48277=>X"00",
48278=>X"00",
48279=>X"00",
48280=>X"00",
48281=>X"00",
48282=>X"00",
48283=>X"00",
48284=>X"00",
48285=>X"00",
48286=>X"00",
48287=>X"00",
48288=>X"00",
48289=>X"00",
48290=>X"00",
48291=>X"00",
48292=>X"00",
48293=>X"00",
48294=>X"00",
48295=>X"00",
48296=>X"00",
48297=>X"00",
48298=>X"00",
48299=>X"00",
48300=>X"00",
48301=>X"00",
48302=>X"00",
48303=>X"00",
48304=>X"00",
48305=>X"00",
48306=>X"00",
48307=>X"00",
48308=>X"00",
48309=>X"00",
48310=>X"00",
48311=>X"00",
48312=>X"00",
48313=>X"00",
48314=>X"00",
48315=>X"00",
48316=>X"00",
48317=>X"00",
48318=>X"00",
48319=>X"00",
48320=>X"00",
48321=>X"00",
48322=>X"00",
48323=>X"00",
48324=>X"00",
48325=>X"00",
48326=>X"00",
48327=>X"00",
48328=>X"00",
48329=>X"00",
48330=>X"00",
48331=>X"00",
48332=>X"00",
48333=>X"00",
48334=>X"00",
48335=>X"00",
48336=>X"00",
48337=>X"00",
48338=>X"00",
48339=>X"00",
48340=>X"00",
48341=>X"00",
48342=>X"00",
48343=>X"00",
48344=>X"00",
48345=>X"00",
48346=>X"00",
48347=>X"00",
48348=>X"00",
48349=>X"00",
48350=>X"00",
48351=>X"00",
48352=>X"00",
48353=>X"00",
48354=>X"00",
48355=>X"00",
48356=>X"00",
48357=>X"00",
48358=>X"00",
48359=>X"00",
48360=>X"00",
48361=>X"00",
48362=>X"00",
48363=>X"00",
48364=>X"00",
48365=>X"00",
48366=>X"00",
48367=>X"00",
48368=>X"00",
48369=>X"00",
48370=>X"00",
48371=>X"00",
48372=>X"00",
48373=>X"00",
48374=>X"00",
48375=>X"00",
48376=>X"00",
48377=>X"00",
48378=>X"00",
48379=>X"00",
48380=>X"00",
48381=>X"00",
48382=>X"00",
48383=>X"00",
48384=>X"00",
48385=>X"00",
48386=>X"00",
48387=>X"00",
48388=>X"00",
48389=>X"00",
48390=>X"00",
48391=>X"00",
48392=>X"00",
48393=>X"00",
48394=>X"00",
48395=>X"00",
48396=>X"00",
48397=>X"00",
48398=>X"00",
48399=>X"00",
48400=>X"00",
48401=>X"00",
48402=>X"00",
48403=>X"00",
48404=>X"00",
48405=>X"00",
48406=>X"00",
48407=>X"00",
48408=>X"00",
48409=>X"00",
48410=>X"00",
48411=>X"00",
48412=>X"00",
48413=>X"00",
48414=>X"00",
48415=>X"00",
48416=>X"00",
48417=>X"00",
48418=>X"00",
48419=>X"00",
48420=>X"00",
48421=>X"00",
48422=>X"00",
48423=>X"00",
48424=>X"00",
48425=>X"00",
48426=>X"00",
48427=>X"00",
48428=>X"00",
48429=>X"00",
48430=>X"00",
48431=>X"00",
48432=>X"00",
48433=>X"00",
48434=>X"00",
48435=>X"00",
48436=>X"00",
48437=>X"00",
48438=>X"00",
48439=>X"00",
48440=>X"00",
48441=>X"00",
48442=>X"00",
48443=>X"00",
48444=>X"00",
48445=>X"00",
48446=>X"00",
48447=>X"00",
48448=>X"00",
48449=>X"00",
48450=>X"00",
48451=>X"00",
48452=>X"00",
48453=>X"00",
48454=>X"00",
48455=>X"00",
48456=>X"00",
48457=>X"00",
48458=>X"00",
48459=>X"00",
48460=>X"00",
48461=>X"00",
48462=>X"00",
48463=>X"00",
48464=>X"00",
48465=>X"00",
48466=>X"00",
48467=>X"00",
48468=>X"00",
48469=>X"00",
48470=>X"00",
48471=>X"00",
48472=>X"00",
48473=>X"00",
48474=>X"00",
48475=>X"00",
48476=>X"00",
48477=>X"00",
48478=>X"00",
48479=>X"00",
48480=>X"00",
48481=>X"00",
48482=>X"00",
48483=>X"00",
48484=>X"00",
48485=>X"00",
48486=>X"00",
48487=>X"00",
48488=>X"00",
48489=>X"00",
48490=>X"00",
48491=>X"00",
48492=>X"00",
48493=>X"00",
48494=>X"00",
48495=>X"00",
48496=>X"00",
48497=>X"00",
48498=>X"00",
48499=>X"00",
48500=>X"00",
48501=>X"00",
48502=>X"00",
48503=>X"00",
48504=>X"00",
48505=>X"00",
48506=>X"00",
48507=>X"00",
48508=>X"00",
48509=>X"00",
48510=>X"00",
48511=>X"00",
48512=>X"00",
48513=>X"00",
48514=>X"00",
48515=>X"00",
48516=>X"00",
48517=>X"00",
48518=>X"00",
48519=>X"00",
48520=>X"00",
48521=>X"00",
48522=>X"00",
48523=>X"00",
48524=>X"00",
48525=>X"00",
48526=>X"00",
48527=>X"00",
48528=>X"00",
48529=>X"00",
48530=>X"00",
48531=>X"00",
48532=>X"00",
48533=>X"00",
48534=>X"00",
48535=>X"00",
48536=>X"00",
48537=>X"00",
48538=>X"00",
48539=>X"00",
48540=>X"00",
48541=>X"00",
48542=>X"00",
48543=>X"00",
48544=>X"00",
48545=>X"00",
48546=>X"00",
48547=>X"00",
48548=>X"00",
48549=>X"00",
48550=>X"00",
48551=>X"00",
48552=>X"00",
48553=>X"00",
48554=>X"00",
48555=>X"00",
48556=>X"00",
48557=>X"00",
48558=>X"00",
48559=>X"00",
48560=>X"00",
48561=>X"00",
48562=>X"00",
48563=>X"00",
48564=>X"00",
48565=>X"00",
48566=>X"00",
48567=>X"00",
48568=>X"00",
48569=>X"00",
48570=>X"00",
48571=>X"00",
48572=>X"00",
48573=>X"00",
48574=>X"00",
48575=>X"00",
48576=>X"00",
48577=>X"00",
48578=>X"00",
48579=>X"00",
48580=>X"00",
48581=>X"00",
48582=>X"00",
48583=>X"00",
48584=>X"00",
48585=>X"00",
48586=>X"00",
48587=>X"00",
48588=>X"00",
48589=>X"00",
48590=>X"00",
48591=>X"00",
48592=>X"00",
48593=>X"00",
48594=>X"00",
48595=>X"00",
48596=>X"00",
48597=>X"00",
48598=>X"00",
48599=>X"00",
48600=>X"00",
48601=>X"00",
48602=>X"00",
48603=>X"00",
48604=>X"00",
48605=>X"00",
48606=>X"00",
48607=>X"00",
48608=>X"00",
48609=>X"00",
48610=>X"00",
48611=>X"00",
48612=>X"00",
48613=>X"00",
48614=>X"00",
48615=>X"00",
48616=>X"00",
48617=>X"00",
48618=>X"00",
48619=>X"00",
48620=>X"00",
48621=>X"00",
48622=>X"00",
48623=>X"00",
48624=>X"00",
48625=>X"00",
48626=>X"00",
48627=>X"00",
48628=>X"00",
48629=>X"00",
48630=>X"00",
48631=>X"00",
48632=>X"00",
48633=>X"00",
48634=>X"00",
48635=>X"00",
48636=>X"00",
48637=>X"00",
48638=>X"00",
48639=>X"00",
48640=>X"00",
48641=>X"00",
48642=>X"00",
48643=>X"00",
48644=>X"00",
48645=>X"00",
48646=>X"00",
48647=>X"00",
48648=>X"00",
48649=>X"00",
48650=>X"00",
48651=>X"00",
48652=>X"00",
48653=>X"00",
48654=>X"00",
48655=>X"00",
48656=>X"00",
48657=>X"00",
48658=>X"00",
48659=>X"00",
48660=>X"00",
48661=>X"00",
48662=>X"00",
48663=>X"00",
48664=>X"00",
48665=>X"00",
48666=>X"00",
48667=>X"00",
48668=>X"00",
48669=>X"00",
48670=>X"00",
48671=>X"00",
48672=>X"00",
48673=>X"00",
48674=>X"00",
48675=>X"00",
48676=>X"00",
48677=>X"00",
48678=>X"00",
48679=>X"00",
48680=>X"00",
48681=>X"00",
48682=>X"00",
48683=>X"00",
48684=>X"00",
48685=>X"00",
48686=>X"00",
48687=>X"00",
48688=>X"00",
48689=>X"00",
48690=>X"00",
48691=>X"00",
48692=>X"00",
48693=>X"00",
48694=>X"00",
48695=>X"00",
48696=>X"00",
48697=>X"00",
48698=>X"00",
48699=>X"00",
48700=>X"00",
48701=>X"00",
48702=>X"00",
48703=>X"00",
48704=>X"00",
48705=>X"00",
48706=>X"00",
48707=>X"00",
48708=>X"00",
48709=>X"00",
48710=>X"00",
48711=>X"00",
48712=>X"00",
48713=>X"00",
48714=>X"00",
48715=>X"00",
48716=>X"00",
48717=>X"00",
48718=>X"00",
48719=>X"00",
48720=>X"00",
48721=>X"00",
48722=>X"00",
48723=>X"00",
48724=>X"00",
48725=>X"00",
48726=>X"00",
48727=>X"00",
48728=>X"00",
48729=>X"00",
48730=>X"00",
48731=>X"00",
48732=>X"00",
48733=>X"00",
48734=>X"00",
48735=>X"00",
48736=>X"00",
48737=>X"00",
48738=>X"00",
48739=>X"00",
48740=>X"00",
48741=>X"00",
48742=>X"00",
48743=>X"00",
48744=>X"00",
48745=>X"00",
48746=>X"00",
48747=>X"00",
48748=>X"00",
48749=>X"00",
48750=>X"00",
48751=>X"00",
48752=>X"00",
48753=>X"00",
48754=>X"00",
48755=>X"00",
48756=>X"00",
48757=>X"00",
48758=>X"00",
48759=>X"00",
48760=>X"00",
48761=>X"00",
48762=>X"00",
48763=>X"00",
48764=>X"00",
48765=>X"00",
48766=>X"00",
48767=>X"00",
48768=>X"00",
48769=>X"00",
48770=>X"00",
48771=>X"00",
48772=>X"00",
48773=>X"00",
48774=>X"00",
48775=>X"00",
48776=>X"00",
48777=>X"00",
48778=>X"00",
48779=>X"00",
48780=>X"00",
48781=>X"00",
48782=>X"00",
48783=>X"00",
48784=>X"00",
48785=>X"00",
48786=>X"00",
48787=>X"00",
48788=>X"00",
48789=>X"00",
48790=>X"00",
48791=>X"00",
48792=>X"00",
48793=>X"00",
48794=>X"00",
48795=>X"00",
48796=>X"00",
48797=>X"00",
48798=>X"00",
48799=>X"00",
48800=>X"00",
48801=>X"00",
48802=>X"00",
48803=>X"00",
48804=>X"00",
48805=>X"00",
48806=>X"00",
48807=>X"00",
48808=>X"00",
48809=>X"00",
48810=>X"00",
48811=>X"00",
48812=>X"00",
48813=>X"00",
48814=>X"00",
48815=>X"00",
48816=>X"00",
48817=>X"00",
48818=>X"00",
48819=>X"00",
48820=>X"00",
48821=>X"00",
48822=>X"00",
48823=>X"00",
48824=>X"00",
48825=>X"00",
48826=>X"00",
48827=>X"00",
48828=>X"00",
48829=>X"00",
48830=>X"00",
48831=>X"00",
48832=>X"00",
48833=>X"00",
48834=>X"00",
48835=>X"00",
48836=>X"00",
48837=>X"00",
48838=>X"00",
48839=>X"00",
48840=>X"00",
48841=>X"00",
48842=>X"00",
48843=>X"00",
48844=>X"00",
48845=>X"00",
48846=>X"00",
48847=>X"00",
48848=>X"00",
48849=>X"00",
48850=>X"00",
48851=>X"00",
48852=>X"00",
48853=>X"00",
48854=>X"00",
48855=>X"00",
48856=>X"00",
48857=>X"00",
48858=>X"00",
48859=>X"00",
48860=>X"00",
48861=>X"00",
48862=>X"00",
48863=>X"00",
48864=>X"00",
48865=>X"00",
48866=>X"00",
48867=>X"00",
48868=>X"00",
48869=>X"00",
48870=>X"00",
48871=>X"00",
48872=>X"00",
48873=>X"00",
48874=>X"00",
48875=>X"00",
48876=>X"00",
48877=>X"00",
48878=>X"00",
48879=>X"00",
48880=>X"00",
48881=>X"00",
48882=>X"00",
48883=>X"00",
48884=>X"00",
48885=>X"00",
48886=>X"00",
48887=>X"00",
48888=>X"00",
48889=>X"00",
48890=>X"00",
48891=>X"00",
48892=>X"00",
48893=>X"00",
48894=>X"00",
48895=>X"00",
48896=>X"00",
48897=>X"00",
48898=>X"00",
48899=>X"00",
48900=>X"00",
48901=>X"00",
48902=>X"00",
48903=>X"00",
48904=>X"00",
48905=>X"00",
48906=>X"00",
48907=>X"00",
48908=>X"00",
48909=>X"00",
48910=>X"00",
48911=>X"00",
48912=>X"00",
48913=>X"00",
48914=>X"00",
48915=>X"00",
48916=>X"00",
48917=>X"00",
48918=>X"00",
48919=>X"00",
48920=>X"00",
48921=>X"00",
48922=>X"00",
48923=>X"00",
48924=>X"00",
48925=>X"00",
48926=>X"00",
48927=>X"00",
48928=>X"00",
48929=>X"00",
48930=>X"00",
48931=>X"00",
48932=>X"00",
48933=>X"00",
48934=>X"00",
48935=>X"00",
48936=>X"00",
48937=>X"00",
48938=>X"00",
48939=>X"00",
48940=>X"00",
48941=>X"00",
48942=>X"00",
48943=>X"00",
48944=>X"00",
48945=>X"00",
48946=>X"00",
48947=>X"00",
48948=>X"00",
48949=>X"00",
48950=>X"00",
48951=>X"00",
48952=>X"00",
48953=>X"00",
48954=>X"00",
48955=>X"00",
48956=>X"00",
48957=>X"00",
48958=>X"00",
48959=>X"00",
48960=>X"00",
48961=>X"00",
48962=>X"00",
48963=>X"00",
48964=>X"00",
48965=>X"00",
48966=>X"00",
48967=>X"00",
48968=>X"00",
48969=>X"00",
48970=>X"00",
48971=>X"00",
48972=>X"00",
48973=>X"00",
48974=>X"00",
48975=>X"00",
48976=>X"00",
48977=>X"00",
48978=>X"00",
48979=>X"00",
48980=>X"00",
48981=>X"00",
48982=>X"00",
48983=>X"00",
48984=>X"00",
48985=>X"00",
48986=>X"00",
48987=>X"00",
48988=>X"00",
48989=>X"00",
48990=>X"00",
48991=>X"00",
48992=>X"00",
48993=>X"00",
48994=>X"00",
48995=>X"00",
48996=>X"00",
48997=>X"00",
48998=>X"00",
48999=>X"00",
49000=>X"00",
49001=>X"00",
49002=>X"00",
49003=>X"00",
49004=>X"00",
49005=>X"00",
49006=>X"00",
49007=>X"00",
49008=>X"00",
49009=>X"00",
49010=>X"00",
49011=>X"00",
49012=>X"00",
49013=>X"00",
49014=>X"00",
49015=>X"00",
49016=>X"00",
49017=>X"00",
49018=>X"00",
49019=>X"00",
49020=>X"00",
49021=>X"00",
49022=>X"00",
49023=>X"00",
49024=>X"00",
49025=>X"00",
49026=>X"00",
49027=>X"00",
49028=>X"00",
49029=>X"00",
49030=>X"00",
49031=>X"00",
49032=>X"00",
49033=>X"00",
49034=>X"00",
49035=>X"00",
49036=>X"00",
49037=>X"00",
49038=>X"00",
49039=>X"00",
49040=>X"00",
49041=>X"00",
49042=>X"00",
49043=>X"00",
49044=>X"00",
49045=>X"00",
49046=>X"00",
49047=>X"00",
49048=>X"00",
49049=>X"00",
49050=>X"00",
49051=>X"00",
49052=>X"00",
49053=>X"00",
49054=>X"00",
49055=>X"00",
49056=>X"00",
49057=>X"00",
49058=>X"00",
49059=>X"00",
49060=>X"00",
49061=>X"00",
49062=>X"00",
49063=>X"00",
49064=>X"00",
49065=>X"00",
49066=>X"00",
49067=>X"00",
49068=>X"00",
49069=>X"00",
49070=>X"00",
49071=>X"00",
49072=>X"00",
49073=>X"00",
49074=>X"00",
49075=>X"00",
49076=>X"00",
49077=>X"00",
49078=>X"00",
49079=>X"00",
49080=>X"00",
49081=>X"00",
49082=>X"00",
49083=>X"00",
49084=>X"00",
49085=>X"00",
49086=>X"00",
49087=>X"00",
49088=>X"00",
49089=>X"00",
49090=>X"00",
49091=>X"00",
49092=>X"00",
49093=>X"00",
49094=>X"00",
49095=>X"00",
49096=>X"00",
49097=>X"00",
49098=>X"00",
49099=>X"00",
49100=>X"00",
49101=>X"00",
49102=>X"00",
49103=>X"00",
49104=>X"00",
49105=>X"00",
49106=>X"00",
49107=>X"00",
49108=>X"00",
49109=>X"00",
49110=>X"00",
49111=>X"00",
49112=>X"00",
49113=>X"00",
49114=>X"00",
49115=>X"00",
49116=>X"00",
49117=>X"00",
49118=>X"00",
49119=>X"00",
49120=>X"00",
49121=>X"00",
49122=>X"00",
49123=>X"00",
49124=>X"00",
49125=>X"00",
49126=>X"00",
49127=>X"00",
49128=>X"00",
49129=>X"00",
49130=>X"00",
49131=>X"00",
49132=>X"00",
49133=>X"00",
49134=>X"00",
49135=>X"00",
49136=>X"00",
49137=>X"00",
49138=>X"00",
49139=>X"00",
49140=>X"00",
49141=>X"00",
49142=>X"00",
49143=>X"00",
49144=>X"00",
49145=>X"00",
49146=>X"00",
49147=>X"00",
49148=>X"00",
49149=>X"00",
49150=>X"00",
49151=>X"00",
49152=>X"00",
49153=>X"00",
49154=>X"00",
49155=>X"00",
49156=>X"00",
49157=>X"00",
49158=>X"00",
49159=>X"00",
49160=>X"00",
49161=>X"00",
49162=>X"00",
49163=>X"00",
49164=>X"00",
49165=>X"00",
49166=>X"00",
49167=>X"00",
49168=>X"00",
49169=>X"00",
49170=>X"00",
49171=>X"00",
49172=>X"00",
49173=>X"00",
49174=>X"00",
49175=>X"00",
49176=>X"00",
49177=>X"00",
49178=>X"00",
49179=>X"00",
49180=>X"00",
49181=>X"00",
49182=>X"00",
49183=>X"00",
49184=>X"00",
49185=>X"00",
49186=>X"00",
49187=>X"00",
49188=>X"00",
49189=>X"00",
49190=>X"00",
49191=>X"00",
49192=>X"00",
49193=>X"00",
49194=>X"00",
49195=>X"00",
49196=>X"00",
49197=>X"00",
49198=>X"00",
49199=>X"00",
49200=>X"00",
49201=>X"00",
49202=>X"00",
49203=>X"00",
49204=>X"00",
49205=>X"00",
49206=>X"00",
49207=>X"00",
49208=>X"00",
49209=>X"00",
49210=>X"00",
49211=>X"00",
49212=>X"00",
49213=>X"00",
49214=>X"00",
49215=>X"00",
49216=>X"00",
49217=>X"00",
49218=>X"00",
49219=>X"00",
49220=>X"00",
49221=>X"00",
49222=>X"00",
49223=>X"00",
49224=>X"00",
49225=>X"00",
49226=>X"00",
49227=>X"00",
49228=>X"00",
49229=>X"00",
49230=>X"00",
49231=>X"00",
49232=>X"00",
49233=>X"00",
49234=>X"00",
49235=>X"00",
49236=>X"00",
49237=>X"00",
49238=>X"00",
49239=>X"00",
49240=>X"00",
49241=>X"00",
49242=>X"00",
49243=>X"00",
49244=>X"00",
49245=>X"00",
49246=>X"00",
49247=>X"00",
49248=>X"00",
49249=>X"00",
49250=>X"00",
49251=>X"00",
49252=>X"00",
49253=>X"00",
49254=>X"00",
49255=>X"00",
49256=>X"00",
49257=>X"00",
49258=>X"00",
49259=>X"00",
49260=>X"00",
49261=>X"00",
49262=>X"00",
49263=>X"00",
49264=>X"00",
49265=>X"00",
49266=>X"00",
49267=>X"00",
49268=>X"00",
49269=>X"00",
49270=>X"00",
49271=>X"00",
49272=>X"00",
49273=>X"00",
49274=>X"00",
49275=>X"00",
49276=>X"00",
49277=>X"00",
49278=>X"00",
49279=>X"00",
49280=>X"00",
49281=>X"00",
49282=>X"00",
49283=>X"00",
49284=>X"00",
49285=>X"00",
49286=>X"00",
49287=>X"00",
49288=>X"00",
49289=>X"00",
49290=>X"00",
49291=>X"00",
49292=>X"00",
49293=>X"00",
49294=>X"00",
49295=>X"00",
49296=>X"00",
49297=>X"00",
49298=>X"00",
49299=>X"00",
49300=>X"00",
49301=>X"00",
49302=>X"00",
49303=>X"00",
49304=>X"00",
49305=>X"00",
49306=>X"00",
49307=>X"00",
49308=>X"00",
49309=>X"00",
49310=>X"00",
49311=>X"00",
49312=>X"00",
49313=>X"00",
49314=>X"00",
49315=>X"00",
49316=>X"00",
49317=>X"00",
49318=>X"00",
49319=>X"00",
49320=>X"00",
49321=>X"00",
49322=>X"00",
49323=>X"00",
49324=>X"00",
49325=>X"00",
49326=>X"00",
49327=>X"00",
49328=>X"00",
49329=>X"00",
49330=>X"00",
49331=>X"00",
49332=>X"00",
49333=>X"00",
49334=>X"00",
49335=>X"00",
49336=>X"00",
49337=>X"00",
49338=>X"00",
49339=>X"00",
49340=>X"00",
49341=>X"00",
49342=>X"00",
49343=>X"00",
49344=>X"00",
49345=>X"00",
49346=>X"00",
49347=>X"00",
49348=>X"00",
49349=>X"00",
49350=>X"00",
49351=>X"00",
49352=>X"00",
49353=>X"00",
49354=>X"00",
49355=>X"00",
49356=>X"00",
49357=>X"00",
49358=>X"00",
49359=>X"00",
49360=>X"00",
49361=>X"00",
49362=>X"00",
49363=>X"00",
49364=>X"00",
49365=>X"00",
49366=>X"00",
49367=>X"00",
49368=>X"00",
49369=>X"00",
49370=>X"00",
49371=>X"00",
49372=>X"00",
49373=>X"00",
49374=>X"00",
49375=>X"00",
49376=>X"00",
49377=>X"00",
49378=>X"00",
49379=>X"00",
49380=>X"00",
49381=>X"00",
49382=>X"00",
49383=>X"00",
49384=>X"00",
49385=>X"00",
49386=>X"00",
49387=>X"00",
49388=>X"00",
49389=>X"00",
49390=>X"00",
49391=>X"00",
49392=>X"00",
49393=>X"00",
49394=>X"00",
49395=>X"00",
49396=>X"00",
49397=>X"00",
49398=>X"00",
49399=>X"00",
49400=>X"00",
49401=>X"00",
49402=>X"00",
49403=>X"00",
49404=>X"00",
49405=>X"00",
49406=>X"00",
49407=>X"00",
49408=>X"00",
49409=>X"00",
49410=>X"00",
49411=>X"00",
49412=>X"00",
49413=>X"00",
49414=>X"00",
49415=>X"00",
49416=>X"00",
49417=>X"00",
49418=>X"00",
49419=>X"00",
49420=>X"00",
49421=>X"00",
49422=>X"00",
49423=>X"00",
49424=>X"00",
49425=>X"00",
49426=>X"00",
49427=>X"00",
49428=>X"00",
49429=>X"00",
49430=>X"00",
49431=>X"00",
49432=>X"00",
49433=>X"00",
49434=>X"00",
49435=>X"00",
49436=>X"00",
49437=>X"00",
49438=>X"00",
49439=>X"00",
49440=>X"00",
49441=>X"00",
49442=>X"00",
49443=>X"00",
49444=>X"00",
49445=>X"00",
49446=>X"00",
49447=>X"00",
49448=>X"00",
49449=>X"00",
49450=>X"00",
49451=>X"00",
49452=>X"00",
49453=>X"00",
49454=>X"00",
49455=>X"00",
49456=>X"00",
49457=>X"00",
49458=>X"00",
49459=>X"00",
49460=>X"00",
49461=>X"00",
49462=>X"00",
49463=>X"00",
49464=>X"00",
49465=>X"00",
49466=>X"00",
49467=>X"00",
49468=>X"00",
49469=>X"00",
49470=>X"00",
49471=>X"00",
49472=>X"00",
49473=>X"00",
49474=>X"00",
49475=>X"00",
49476=>X"00",
49477=>X"00",
49478=>X"00",
49479=>X"00",
49480=>X"00",
49481=>X"00",
49482=>X"00",
49483=>X"00",
49484=>X"00",
49485=>X"00",
49486=>X"00",
49487=>X"00",
49488=>X"00",
49489=>X"00",
49490=>X"00",
49491=>X"00",
49492=>X"00",
49493=>X"00",
49494=>X"00",
49495=>X"00",
49496=>X"00",
49497=>X"00",
49498=>X"00",
49499=>X"00",
49500=>X"00",
49501=>X"00",
49502=>X"00",
49503=>X"00",
49504=>X"00",
49505=>X"00",
49506=>X"00",
49507=>X"00",
49508=>X"00",
49509=>X"00",
49510=>X"00",
49511=>X"00",
49512=>X"00",
49513=>X"00",
49514=>X"00",
49515=>X"00",
49516=>X"00",
49517=>X"00",
49518=>X"00",
49519=>X"00",
49520=>X"00",
49521=>X"00",
49522=>X"00",
49523=>X"00",
49524=>X"00",
49525=>X"00",
49526=>X"00",
49527=>X"00",
49528=>X"00",
49529=>X"00",
49530=>X"00",
49531=>X"00",
49532=>X"00",
49533=>X"00",
49534=>X"00",
49535=>X"00",
49536=>X"00",
49537=>X"00",
49538=>X"00",
49539=>X"00",
49540=>X"00",
49541=>X"00",
49542=>X"00",
49543=>X"00",
49544=>X"00",
49545=>X"00",
49546=>X"00",
49547=>X"00",
49548=>X"00",
49549=>X"00",
49550=>X"00",
49551=>X"00",
49552=>X"00",
49553=>X"00",
49554=>X"00",
49555=>X"00",
49556=>X"00",
49557=>X"00",
49558=>X"00",
49559=>X"00",
49560=>X"00",
49561=>X"00",
49562=>X"00",
49563=>X"00",
49564=>X"00",
49565=>X"00",
49566=>X"00",
49567=>X"00",
49568=>X"00",
49569=>X"00",
49570=>X"00",
49571=>X"00",
49572=>X"00",
49573=>X"00",
49574=>X"00",
49575=>X"00",
49576=>X"00",
49577=>X"00",
49578=>X"00",
49579=>X"00",
49580=>X"00",
49581=>X"00",
49582=>X"00",
49583=>X"00",
49584=>X"00",
49585=>X"00",
49586=>X"00",
49587=>X"00",
49588=>X"00",
49589=>X"00",
49590=>X"00",
49591=>X"00",
49592=>X"00",
49593=>X"00",
49594=>X"00",
49595=>X"00",
49596=>X"00",
49597=>X"00",
49598=>X"00",
49599=>X"00",
49600=>X"00",
49601=>X"00",
49602=>X"00",
49603=>X"00",
49604=>X"00",
49605=>X"00",
49606=>X"00",
49607=>X"00",
49608=>X"00",
49609=>X"00",
49610=>X"00",
49611=>X"00",
49612=>X"00",
49613=>X"00",
49614=>X"00",
49615=>X"00",
49616=>X"00",
49617=>X"00",
49618=>X"00",
49619=>X"00",
49620=>X"00",
49621=>X"00",
49622=>X"00",
49623=>X"00",
49624=>X"00",
49625=>X"00",
49626=>X"00",
49627=>X"00",
49628=>X"00",
49629=>X"00",
49630=>X"00",
49631=>X"00",
49632=>X"00",
49633=>X"00",
49634=>X"00",
49635=>X"00",
49636=>X"00",
49637=>X"00",
49638=>X"00",
49639=>X"00",
49640=>X"00",
49641=>X"00",
49642=>X"00",
49643=>X"00",
49644=>X"00",
49645=>X"00",
49646=>X"00",
49647=>X"00",
49648=>X"00",
49649=>X"00",
49650=>X"00",
49651=>X"00",
49652=>X"00",
49653=>X"00",
49654=>X"00",
49655=>X"00",
49656=>X"00",
49657=>X"00",
49658=>X"00",
49659=>X"00",
49660=>X"00",
49661=>X"00",
49662=>X"00",
49663=>X"00",
49664=>X"00",
49665=>X"00",
49666=>X"00",
49667=>X"00",
49668=>X"00",
49669=>X"00",
49670=>X"00",
49671=>X"00",
49672=>X"00",
49673=>X"00",
49674=>X"00",
49675=>X"00",
49676=>X"00",
49677=>X"00",
49678=>X"00",
49679=>X"00",
49680=>X"00",
49681=>X"00",
49682=>X"00",
49683=>X"00",
49684=>X"00",
49685=>X"00",
49686=>X"00",
49687=>X"00",
49688=>X"00",
49689=>X"00",
49690=>X"00",
49691=>X"00",
49692=>X"00",
49693=>X"00",
49694=>X"00",
49695=>X"00",
49696=>X"00",
49697=>X"00",
49698=>X"00",
49699=>X"00",
49700=>X"00",
49701=>X"00",
49702=>X"00",
49703=>X"00",
49704=>X"00",
49705=>X"00",
49706=>X"00",
49707=>X"00",
49708=>X"00",
49709=>X"00",
49710=>X"00",
49711=>X"00",
49712=>X"00",
49713=>X"00",
49714=>X"00",
49715=>X"00",
49716=>X"00",
49717=>X"00",
49718=>X"00",
49719=>X"00",
49720=>X"00",
49721=>X"00",
49722=>X"00",
49723=>X"00",
49724=>X"00",
49725=>X"00",
49726=>X"00",
49727=>X"00",
49728=>X"00",
49729=>X"00",
49730=>X"00",
49731=>X"00",
49732=>X"00",
49733=>X"00",
49734=>X"00",
49735=>X"00",
49736=>X"00",
49737=>X"00",
49738=>X"00",
49739=>X"00",
49740=>X"00",
49741=>X"00",
49742=>X"00",
49743=>X"00",
49744=>X"00",
49745=>X"00",
49746=>X"00",
49747=>X"00",
49748=>X"00",
49749=>X"00",
49750=>X"00",
49751=>X"00",
49752=>X"00",
49753=>X"00",
49754=>X"00",
49755=>X"00",
49756=>X"00",
49757=>X"00",
49758=>X"00",
49759=>X"00",
49760=>X"00",
49761=>X"00",
49762=>X"00",
49763=>X"00",
49764=>X"00",
49765=>X"00",
49766=>X"00",
49767=>X"00",
49768=>X"00",
49769=>X"00",
49770=>X"00",
49771=>X"00",
49772=>X"00",
49773=>X"00",
49774=>X"00",
49775=>X"00",
49776=>X"00",
49777=>X"00",
49778=>X"00",
49779=>X"00",
49780=>X"00",
49781=>X"00",
49782=>X"00",
49783=>X"00",
49784=>X"00",
49785=>X"00",
49786=>X"00",
49787=>X"00",
49788=>X"00",
49789=>X"00",
49790=>X"00",
49791=>X"00",
49792=>X"00",
49793=>X"00",
49794=>X"00",
49795=>X"00",
49796=>X"00",
49797=>X"00",
49798=>X"00",
49799=>X"00",
49800=>X"00",
49801=>X"00",
49802=>X"00",
49803=>X"00",
49804=>X"00",
49805=>X"00",
49806=>X"00",
49807=>X"00",
49808=>X"00",
49809=>X"00",
49810=>X"00",
49811=>X"00",
49812=>X"00",
49813=>X"00",
49814=>X"00",
49815=>X"00",
49816=>X"00",
49817=>X"00",
49818=>X"00",
49819=>X"00",
49820=>X"00",
49821=>X"00",
49822=>X"00",
49823=>X"00",
49824=>X"00",
49825=>X"00",
49826=>X"00",
49827=>X"00",
49828=>X"00",
49829=>X"00",
49830=>X"00",
49831=>X"00",
49832=>X"00",
49833=>X"00",
49834=>X"00",
49835=>X"00",
49836=>X"00",
49837=>X"00",
49838=>X"00",
49839=>X"00",
49840=>X"00",
49841=>X"00",
49842=>X"00",
49843=>X"00",
49844=>X"00",
49845=>X"00",
49846=>X"00",
49847=>X"00",
49848=>X"00",
49849=>X"00",
49850=>X"00",
49851=>X"00",
49852=>X"00",
49853=>X"00",
49854=>X"00",
49855=>X"00",
49856=>X"00",
49857=>X"00",
49858=>X"00",
49859=>X"00",
49860=>X"00",
49861=>X"00",
49862=>X"00",
49863=>X"00",
49864=>X"00",
49865=>X"00",
49866=>X"00",
49867=>X"00",
49868=>X"00",
49869=>X"00",
49870=>X"00",
49871=>X"00",
49872=>X"00",
49873=>X"00",
49874=>X"00",
49875=>X"00",
49876=>X"00",
49877=>X"00",
49878=>X"00",
49879=>X"00",
49880=>X"00",
49881=>X"00",
49882=>X"00",
49883=>X"00",
49884=>X"00",
49885=>X"00",
49886=>X"00",
49887=>X"00",
49888=>X"00",
49889=>X"00",
49890=>X"00",
49891=>X"00",
49892=>X"00",
49893=>X"00",
49894=>X"00",
49895=>X"00",
49896=>X"00",
49897=>X"00",
49898=>X"00",
49899=>X"00",
49900=>X"00",
49901=>X"00",
49902=>X"00",
49903=>X"00",
49904=>X"00",
49905=>X"00",
49906=>X"00",
49907=>X"00",
49908=>X"00",
49909=>X"00",
49910=>X"00",
49911=>X"00",
49912=>X"00",
49913=>X"00",
49914=>X"00",
49915=>X"00",
49916=>X"00",
49917=>X"00",
49918=>X"00",
49919=>X"00",
49920=>X"00",
49921=>X"00",
49922=>X"00",
49923=>X"00",
49924=>X"00",
49925=>X"00",
49926=>X"00",
49927=>X"00",
49928=>X"00",
49929=>X"00",
49930=>X"00",
49931=>X"00",
49932=>X"00",
49933=>X"00",
49934=>X"00",
49935=>X"00",
49936=>X"00",
49937=>X"00",
49938=>X"00",
49939=>X"00",
49940=>X"00",
49941=>X"00",
49942=>X"00",
49943=>X"00",
49944=>X"00",
49945=>X"00",
49946=>X"00",
49947=>X"00",
49948=>X"00",
49949=>X"00",
49950=>X"00",
49951=>X"00",
49952=>X"00",
49953=>X"00",
49954=>X"00",
49955=>X"00",
49956=>X"00",
49957=>X"00",
49958=>X"00",
49959=>X"00",
49960=>X"00",
49961=>X"00",
49962=>X"00",
49963=>X"00",
49964=>X"00",
49965=>X"00",
49966=>X"00",
49967=>X"00",
49968=>X"00",
49969=>X"00",
49970=>X"00",
49971=>X"00",
49972=>X"00",
49973=>X"00",
49974=>X"00",
49975=>X"00",
49976=>X"00",
49977=>X"00",
49978=>X"00",
49979=>X"00",
49980=>X"00",
49981=>X"00",
49982=>X"00",
49983=>X"00",
49984=>X"00",
49985=>X"00",
49986=>X"00",
49987=>X"00",
49988=>X"00",
49989=>X"00",
49990=>X"00",
49991=>X"00",
49992=>X"00",
49993=>X"00",
49994=>X"00",
49995=>X"00",
49996=>X"00",
49997=>X"00",
49998=>X"00",
49999=>X"00",
50000=>X"00",
50001=>X"00",
50002=>X"00",
50003=>X"00",
50004=>X"00",
50005=>X"00",
50006=>X"00",
50007=>X"00",
50008=>X"00",
50009=>X"00",
50010=>X"00",
50011=>X"00",
50012=>X"00",
50013=>X"00",
50014=>X"00",
50015=>X"00",
50016=>X"00",
50017=>X"00",
50018=>X"00",
50019=>X"00",
50020=>X"00",
50021=>X"00",
50022=>X"00",
50023=>X"00",
50024=>X"00",
50025=>X"00",
50026=>X"00",
50027=>X"00",
50028=>X"00",
50029=>X"00",
50030=>X"00",
50031=>X"00",
50032=>X"00",
50033=>X"00",
50034=>X"00",
50035=>X"00",
50036=>X"00",
50037=>X"00",
50038=>X"00",
50039=>X"00",
50040=>X"00",
50041=>X"00",
50042=>X"00",
50043=>X"00",
50044=>X"00",
50045=>X"00",
50046=>X"00",
50047=>X"00",
50048=>X"00",
50049=>X"00",
50050=>X"00",
50051=>X"00",
50052=>X"00",
50053=>X"00",
50054=>X"00",
50055=>X"00",
50056=>X"00",
50057=>X"00",
50058=>X"00",
50059=>X"00",
50060=>X"00",
50061=>X"00",
50062=>X"00",
50063=>X"00",
50064=>X"00",
50065=>X"00",
50066=>X"00",
50067=>X"00",
50068=>X"00",
50069=>X"00",
50070=>X"00",
50071=>X"00",
50072=>X"00",
50073=>X"00",
50074=>X"00",
50075=>X"00",
50076=>X"00",
50077=>X"00",
50078=>X"00",
50079=>X"00",
50080=>X"00",
50081=>X"00",
50082=>X"00",
50083=>X"00",
50084=>X"00",
50085=>X"00",
50086=>X"00",
50087=>X"00",
50088=>X"00",
50089=>X"00",
50090=>X"00",
50091=>X"00",
50092=>X"00",
50093=>X"00",
50094=>X"00",
50095=>X"00",
50096=>X"00",
50097=>X"00",
50098=>X"00",
50099=>X"00",
50100=>X"00",
50101=>X"00",
50102=>X"00",
50103=>X"00",
50104=>X"00",
50105=>X"00",
50106=>X"00",
50107=>X"00",
50108=>X"00",
50109=>X"00",
50110=>X"00",
50111=>X"00",
50112=>X"00",
50113=>X"00",
50114=>X"00",
50115=>X"00",
50116=>X"00",
50117=>X"00",
50118=>X"00",
50119=>X"00",
50120=>X"00",
50121=>X"00",
50122=>X"00",
50123=>X"00",
50124=>X"00",
50125=>X"00",
50126=>X"00",
50127=>X"00",
50128=>X"00",
50129=>X"00",
50130=>X"00",
50131=>X"00",
50132=>X"00",
50133=>X"00",
50134=>X"00",
50135=>X"00",
50136=>X"00",
50137=>X"00",
50138=>X"00",
50139=>X"00",
50140=>X"00",
50141=>X"00",
50142=>X"00",
50143=>X"00",
50144=>X"00",
50145=>X"00",
50146=>X"00",
50147=>X"00",
50148=>X"00",
50149=>X"00",
50150=>X"00",
50151=>X"00",
50152=>X"00",
50153=>X"00",
50154=>X"00",
50155=>X"00",
50156=>X"00",
50157=>X"00",
50158=>X"00",
50159=>X"00",
50160=>X"00",
50161=>X"00",
50162=>X"00",
50163=>X"00",
50164=>X"00",
50165=>X"00",
50166=>X"00",
50167=>X"00",
50168=>X"00",
50169=>X"00",
50170=>X"00",
50171=>X"00",
50172=>X"00",
50173=>X"00",
50174=>X"00",
50175=>X"00",
50176=>X"00",
50177=>X"00",
50178=>X"00",
50179=>X"00",
50180=>X"00",
50181=>X"00",
50182=>X"00",
50183=>X"00",
50184=>X"00",
50185=>X"00",
50186=>X"00",
50187=>X"00",
50188=>X"00",
50189=>X"00",
50190=>X"00",
50191=>X"00",
50192=>X"00",
50193=>X"00",
50194=>X"00",
50195=>X"00",
50196=>X"00",
50197=>X"00",
50198=>X"00",
50199=>X"00",
50200=>X"00",
50201=>X"00",
50202=>X"00",
50203=>X"00",
50204=>X"00",
50205=>X"00",
50206=>X"00",
50207=>X"00",
50208=>X"00",
50209=>X"00",
50210=>X"00",
50211=>X"00",
50212=>X"00",
50213=>X"00",
50214=>X"00",
50215=>X"00",
50216=>X"00",
50217=>X"00",
50218=>X"00",
50219=>X"00",
50220=>X"00",
50221=>X"00",
50222=>X"00",
50223=>X"00",
50224=>X"00",
50225=>X"00",
50226=>X"00",
50227=>X"00",
50228=>X"00",
50229=>X"00",
50230=>X"00",
50231=>X"00",
50232=>X"00",
50233=>X"00",
50234=>X"00",
50235=>X"00",
50236=>X"00",
50237=>X"00",
50238=>X"00",
50239=>X"00",
50240=>X"00",
50241=>X"00",
50242=>X"00",
50243=>X"00",
50244=>X"00",
50245=>X"00",
50246=>X"00",
50247=>X"00",
50248=>X"00",
50249=>X"00",
50250=>X"00",
50251=>X"00",
50252=>X"00",
50253=>X"00",
50254=>X"00",
50255=>X"00",
50256=>X"00",
50257=>X"00",
50258=>X"00",
50259=>X"00",
50260=>X"00",
50261=>X"00",
50262=>X"00",
50263=>X"00",
50264=>X"00",
50265=>X"00",
50266=>X"00",
50267=>X"00",
50268=>X"00",
50269=>X"00",
50270=>X"00",
50271=>X"00",
50272=>X"00",
50273=>X"00",
50274=>X"00",
50275=>X"00",
50276=>X"00",
50277=>X"00",
50278=>X"00",
50279=>X"00",
50280=>X"00",
50281=>X"00",
50282=>X"00",
50283=>X"00",
50284=>X"00",
50285=>X"00",
50286=>X"00",
50287=>X"00",
50288=>X"00",
50289=>X"00",
50290=>X"00",
50291=>X"00",
50292=>X"00",
50293=>X"00",
50294=>X"00",
50295=>X"00",
50296=>X"00",
50297=>X"00",
50298=>X"00",
50299=>X"00",
50300=>X"00",
50301=>X"00",
50302=>X"00",
50303=>X"00",
50304=>X"00",
50305=>X"00",
50306=>X"00",
50307=>X"00",
50308=>X"00",
50309=>X"00",
50310=>X"00",
50311=>X"00",
50312=>X"00",
50313=>X"00",
50314=>X"00",
50315=>X"00",
50316=>X"00",
50317=>X"00",
50318=>X"00",
50319=>X"00",
50320=>X"00",
50321=>X"00",
50322=>X"00",
50323=>X"00",
50324=>X"00",
50325=>X"00",
50326=>X"00",
50327=>X"00",
50328=>X"00",
50329=>X"00",
50330=>X"00",
50331=>X"00",
50332=>X"00",
50333=>X"00",
50334=>X"00",
50335=>X"00",
50336=>X"00",
50337=>X"00",
50338=>X"00",
50339=>X"00",
50340=>X"00",
50341=>X"00",
50342=>X"00",
50343=>X"00",
50344=>X"00",
50345=>X"00",
50346=>X"00",
50347=>X"00",
50348=>X"00",
50349=>X"00",
50350=>X"00",
50351=>X"00",
50352=>X"00",
50353=>X"00",
50354=>X"00",
50355=>X"00",
50356=>X"00",
50357=>X"00",
50358=>X"00",
50359=>X"00",
50360=>X"00",
50361=>X"00",
50362=>X"00",
50363=>X"00",
50364=>X"00",
50365=>X"00",
50366=>X"00",
50367=>X"00",
50368=>X"00",
50369=>X"00",
50370=>X"00",
50371=>X"00",
50372=>X"00",
50373=>X"00",
50374=>X"00",
50375=>X"00",
50376=>X"00",
50377=>X"00",
50378=>X"00",
50379=>X"00",
50380=>X"00",
50381=>X"00",
50382=>X"00",
50383=>X"00",
50384=>X"00",
50385=>X"00",
50386=>X"00",
50387=>X"00",
50388=>X"00",
50389=>X"00",
50390=>X"00",
50391=>X"00",
50392=>X"00",
50393=>X"00",
50394=>X"00",
50395=>X"00",
50396=>X"00",
50397=>X"00",
50398=>X"00",
50399=>X"00",
50400=>X"00",
50401=>X"00",
50402=>X"00",
50403=>X"00",
50404=>X"00",
50405=>X"00",
50406=>X"00",
50407=>X"00",
50408=>X"00",
50409=>X"00",
50410=>X"00",
50411=>X"00",
50412=>X"00",
50413=>X"00",
50414=>X"00",
50415=>X"00",
50416=>X"00",
50417=>X"00",
50418=>X"00",
50419=>X"00",
50420=>X"00",
50421=>X"00",
50422=>X"00",
50423=>X"00",
50424=>X"00",
50425=>X"00",
50426=>X"00",
50427=>X"00",
50428=>X"00",
50429=>X"00",
50430=>X"00",
50431=>X"00",
50432=>X"00",
50433=>X"00",
50434=>X"00",
50435=>X"00",
50436=>X"00",
50437=>X"00",
50438=>X"00",
50439=>X"00",
50440=>X"00",
50441=>X"00",
50442=>X"00",
50443=>X"00",
50444=>X"00",
50445=>X"00",
50446=>X"00",
50447=>X"00",
50448=>X"00",
50449=>X"00",
50450=>X"00",
50451=>X"00",
50452=>X"00",
50453=>X"00",
50454=>X"00",
50455=>X"00",
50456=>X"00",
50457=>X"00",
50458=>X"00",
50459=>X"00",
50460=>X"00",
50461=>X"00",
50462=>X"00",
50463=>X"00",
50464=>X"00",
50465=>X"00",
50466=>X"00",
50467=>X"00",
50468=>X"00",
50469=>X"00",
50470=>X"00",
50471=>X"00",
50472=>X"00",
50473=>X"00",
50474=>X"00",
50475=>X"00",
50476=>X"00",
50477=>X"00",
50478=>X"00",
50479=>X"00",
50480=>X"00",
50481=>X"00",
50482=>X"00",
50483=>X"00",
50484=>X"00",
50485=>X"00",
50486=>X"00",
50487=>X"00",
50488=>X"00",
50489=>X"00",
50490=>X"00",
50491=>X"00",
50492=>X"00",
50493=>X"00",
50494=>X"00",
50495=>X"00",
50496=>X"00",
50497=>X"00",
50498=>X"00",
50499=>X"00",
50500=>X"00",
50501=>X"00",
50502=>X"00",
50503=>X"00",
50504=>X"00",
50505=>X"00",
50506=>X"00",
50507=>X"00",
50508=>X"00",
50509=>X"00",
50510=>X"00",
50511=>X"00",
50512=>X"00",
50513=>X"00",
50514=>X"00",
50515=>X"00",
50516=>X"00",
50517=>X"00",
50518=>X"00",
50519=>X"00",
50520=>X"00",
50521=>X"00",
50522=>X"00",
50523=>X"00",
50524=>X"00",
50525=>X"00",
50526=>X"00",
50527=>X"00",
50528=>X"00",
50529=>X"00",
50530=>X"00",
50531=>X"00",
50532=>X"00",
50533=>X"00",
50534=>X"00",
50535=>X"00",
50536=>X"00",
50537=>X"00",
50538=>X"00",
50539=>X"00",
50540=>X"00",
50541=>X"00",
50542=>X"00",
50543=>X"00",
50544=>X"00",
50545=>X"00",
50546=>X"00",
50547=>X"00",
50548=>X"00",
50549=>X"00",
50550=>X"00",
50551=>X"00",
50552=>X"00",
50553=>X"00",
50554=>X"00",
50555=>X"00",
50556=>X"00",
50557=>X"00",
50558=>X"00",
50559=>X"00",
50560=>X"00",
50561=>X"00",
50562=>X"00",
50563=>X"00",
50564=>X"00",
50565=>X"00",
50566=>X"00",
50567=>X"00",
50568=>X"00",
50569=>X"00",
50570=>X"00",
50571=>X"00",
50572=>X"00",
50573=>X"00",
50574=>X"00",
50575=>X"00",
50576=>X"00",
50577=>X"00",
50578=>X"00",
50579=>X"00",
50580=>X"00",
50581=>X"00",
50582=>X"00",
50583=>X"00",
50584=>X"00",
50585=>X"00",
50586=>X"00",
50587=>X"00",
50588=>X"00",
50589=>X"00",
50590=>X"00",
50591=>X"00",
50592=>X"00",
50593=>X"00",
50594=>X"00",
50595=>X"00",
50596=>X"00",
50597=>X"00",
50598=>X"00",
50599=>X"00",
50600=>X"00",
50601=>X"00",
50602=>X"00",
50603=>X"00",
50604=>X"00",
50605=>X"00",
50606=>X"00",
50607=>X"00",
50608=>X"00",
50609=>X"00",
50610=>X"00",
50611=>X"00",
50612=>X"00",
50613=>X"00",
50614=>X"00",
50615=>X"00",
50616=>X"00",
50617=>X"00",
50618=>X"00",
50619=>X"00",
50620=>X"00",
50621=>X"00",
50622=>X"00",
50623=>X"00",
50624=>X"00",
50625=>X"00",
50626=>X"00",
50627=>X"00",
50628=>X"00",
50629=>X"00",
50630=>X"00",
50631=>X"00",
50632=>X"00",
50633=>X"00",
50634=>X"00",
50635=>X"00",
50636=>X"00",
50637=>X"00",
50638=>X"00",
50639=>X"00",
50640=>X"00",
50641=>X"00",
50642=>X"00",
50643=>X"00",
50644=>X"00",
50645=>X"00",
50646=>X"00",
50647=>X"00",
50648=>X"00",
50649=>X"00",
50650=>X"00",
50651=>X"00",
50652=>X"00",
50653=>X"00",
50654=>X"00",
50655=>X"00",
50656=>X"00",
50657=>X"00",
50658=>X"00",
50659=>X"00",
50660=>X"00",
50661=>X"00",
50662=>X"00",
50663=>X"00",
50664=>X"00",
50665=>X"00",
50666=>X"00",
50667=>X"00",
50668=>X"00",
50669=>X"00",
50670=>X"00",
50671=>X"00",
50672=>X"00",
50673=>X"00",
50674=>X"00",
50675=>X"00",
50676=>X"00",
50677=>X"00",
50678=>X"00",
50679=>X"00",
50680=>X"00",
50681=>X"00",
50682=>X"00",
50683=>X"00",
50684=>X"00",
50685=>X"00",
50686=>X"00",
50687=>X"00",
50688=>X"00",
50689=>X"00",
50690=>X"00",
50691=>X"00",
50692=>X"00",
50693=>X"00",
50694=>X"00",
50695=>X"00",
50696=>X"00",
50697=>X"00",
50698=>X"00",
50699=>X"00",
50700=>X"00",
50701=>X"00",
50702=>X"00",
50703=>X"00",
50704=>X"00",
50705=>X"00",
50706=>X"00",
50707=>X"00",
50708=>X"00",
50709=>X"00",
50710=>X"00",
50711=>X"00",
50712=>X"00",
50713=>X"00",
50714=>X"00",
50715=>X"00",
50716=>X"00",
50717=>X"00",
50718=>X"00",
50719=>X"00",
50720=>X"00",
50721=>X"00",
50722=>X"00",
50723=>X"00",
50724=>X"00",
50725=>X"00",
50726=>X"00",
50727=>X"00",
50728=>X"00",
50729=>X"00",
50730=>X"00",
50731=>X"00",
50732=>X"00",
50733=>X"00",
50734=>X"00",
50735=>X"00",
50736=>X"00",
50737=>X"00",
50738=>X"00",
50739=>X"00",
50740=>X"00",
50741=>X"00",
50742=>X"00",
50743=>X"00",
50744=>X"00",
50745=>X"00",
50746=>X"00",
50747=>X"00",
50748=>X"00",
50749=>X"00",
50750=>X"00",
50751=>X"00",
50752=>X"00",
50753=>X"00",
50754=>X"00",
50755=>X"00",
50756=>X"00",
50757=>X"00",
50758=>X"00",
50759=>X"00",
50760=>X"00",
50761=>X"00",
50762=>X"00",
50763=>X"00",
50764=>X"00",
50765=>X"00",
50766=>X"00",
50767=>X"00",
50768=>X"00",
50769=>X"00",
50770=>X"00",
50771=>X"00",
50772=>X"00",
50773=>X"00",
50774=>X"00",
50775=>X"00",
50776=>X"00",
50777=>X"00",
50778=>X"00",
50779=>X"00",
50780=>X"00",
50781=>X"00",
50782=>X"00",
50783=>X"00",
50784=>X"00",
50785=>X"00",
50786=>X"00",
50787=>X"00",
50788=>X"00",
50789=>X"00",
50790=>X"00",
50791=>X"00",
50792=>X"00",
50793=>X"00",
50794=>X"00",
50795=>X"00",
50796=>X"00",
50797=>X"00",
50798=>X"00",
50799=>X"00",
50800=>X"00",
50801=>X"00",
50802=>X"00",
50803=>X"00",
50804=>X"00",
50805=>X"00",
50806=>X"00",
50807=>X"00",
50808=>X"00",
50809=>X"00",
50810=>X"00",
50811=>X"00",
50812=>X"00",
50813=>X"00",
50814=>X"00",
50815=>X"00",
50816=>X"00",
50817=>X"00",
50818=>X"00",
50819=>X"00",
50820=>X"00",
50821=>X"00",
50822=>X"00",
50823=>X"00",
50824=>X"00",
50825=>X"00",
50826=>X"00",
50827=>X"00",
50828=>X"00",
50829=>X"00",
50830=>X"00",
50831=>X"00",
50832=>X"00",
50833=>X"00",
50834=>X"00",
50835=>X"00",
50836=>X"00",
50837=>X"00",
50838=>X"00",
50839=>X"00",
50840=>X"00",
50841=>X"00",
50842=>X"00",
50843=>X"00",
50844=>X"00",
50845=>X"00",
50846=>X"00",
50847=>X"00",
50848=>X"00",
50849=>X"00",
50850=>X"00",
50851=>X"00",
50852=>X"00",
50853=>X"00",
50854=>X"00",
50855=>X"00",
50856=>X"00",
50857=>X"00",
50858=>X"00",
50859=>X"00",
50860=>X"00",
50861=>X"00",
50862=>X"00",
50863=>X"00",
50864=>X"00",
50865=>X"00",
50866=>X"00",
50867=>X"00",
50868=>X"00",
50869=>X"00",
50870=>X"00",
50871=>X"00",
50872=>X"00",
50873=>X"00",
50874=>X"00",
50875=>X"00",
50876=>X"00",
50877=>X"00",
50878=>X"00",
50879=>X"00",
50880=>X"00",
50881=>X"00",
50882=>X"00",
50883=>X"00",
50884=>X"00",
50885=>X"00",
50886=>X"00",
50887=>X"00",
50888=>X"00",
50889=>X"00",
50890=>X"00",
50891=>X"00",
50892=>X"00",
50893=>X"00",
50894=>X"00",
50895=>X"00",
50896=>X"00",
50897=>X"00",
50898=>X"00",
50899=>X"00",
50900=>X"00",
50901=>X"00",
50902=>X"00",
50903=>X"00",
50904=>X"00",
50905=>X"00",
50906=>X"00",
50907=>X"00",
50908=>X"00",
50909=>X"00",
50910=>X"00",
50911=>X"00",
50912=>X"00",
50913=>X"00",
50914=>X"00",
50915=>X"00",
50916=>X"00",
50917=>X"00",
50918=>X"00",
50919=>X"00",
50920=>X"00",
50921=>X"00",
50922=>X"00",
50923=>X"00",
50924=>X"00",
50925=>X"00",
50926=>X"00",
50927=>X"00",
50928=>X"00",
50929=>X"00",
50930=>X"00",
50931=>X"00",
50932=>X"00",
50933=>X"00",
50934=>X"00",
50935=>X"00",
50936=>X"00",
50937=>X"00",
50938=>X"00",
50939=>X"00",
50940=>X"00",
50941=>X"00",
50942=>X"00",
50943=>X"00",
50944=>X"00",
50945=>X"00",
50946=>X"00",
50947=>X"00",
50948=>X"00",
50949=>X"00",
50950=>X"00",
50951=>X"00",
50952=>X"00",
50953=>X"00",
50954=>X"00",
50955=>X"00",
50956=>X"00",
50957=>X"00",
50958=>X"00",
50959=>X"00",
50960=>X"00",
50961=>X"00",
50962=>X"00",
50963=>X"00",
50964=>X"00",
50965=>X"00",
50966=>X"00",
50967=>X"00",
50968=>X"00",
50969=>X"00",
50970=>X"00",
50971=>X"00",
50972=>X"00",
50973=>X"00",
50974=>X"00",
50975=>X"00",
50976=>X"00",
50977=>X"00",
50978=>X"00",
50979=>X"00",
50980=>X"00",
50981=>X"00",
50982=>X"00",
50983=>X"00",
50984=>X"00",
50985=>X"00",
50986=>X"00",
50987=>X"00",
50988=>X"00",
50989=>X"00",
50990=>X"00",
50991=>X"00",
50992=>X"00",
50993=>X"00",
50994=>X"00",
50995=>X"00",
50996=>X"00",
50997=>X"00",
50998=>X"00",
50999=>X"00",
51000=>X"00",
51001=>X"00",
51002=>X"00",
51003=>X"00",
51004=>X"00",
51005=>X"00",
51006=>X"00",
51007=>X"00",
51008=>X"00",
51009=>X"00",
51010=>X"00",
51011=>X"00",
51012=>X"00",
51013=>X"00",
51014=>X"00",
51015=>X"00",
51016=>X"00",
51017=>X"00",
51018=>X"00",
51019=>X"00",
51020=>X"00",
51021=>X"00",
51022=>X"00",
51023=>X"00",
51024=>X"00",
51025=>X"00",
51026=>X"00",
51027=>X"00",
51028=>X"00",
51029=>X"00",
51030=>X"00",
51031=>X"00",
51032=>X"00",
51033=>X"00",
51034=>X"00",
51035=>X"00",
51036=>X"00",
51037=>X"00",
51038=>X"00",
51039=>X"00",
51040=>X"00",
51041=>X"00",
51042=>X"00",
51043=>X"00",
51044=>X"00",
51045=>X"00",
51046=>X"00",
51047=>X"00",
51048=>X"00",
51049=>X"00",
51050=>X"00",
51051=>X"00",
51052=>X"00",
51053=>X"00",
51054=>X"00",
51055=>X"00",
51056=>X"00",
51057=>X"00",
51058=>X"00",
51059=>X"00",
51060=>X"00",
51061=>X"00",
51062=>X"00",
51063=>X"00",
51064=>X"00",
51065=>X"00",
51066=>X"00",
51067=>X"00",
51068=>X"00",
51069=>X"00",
51070=>X"00",
51071=>X"00",
51072=>X"00",
51073=>X"00",
51074=>X"00",
51075=>X"00",
51076=>X"00",
51077=>X"00",
51078=>X"00",
51079=>X"00",
51080=>X"00",
51081=>X"00",
51082=>X"00",
51083=>X"00",
51084=>X"00",
51085=>X"00",
51086=>X"00",
51087=>X"00",
51088=>X"00",
51089=>X"00",
51090=>X"00",
51091=>X"00",
51092=>X"00",
51093=>X"00",
51094=>X"00",
51095=>X"00",
51096=>X"00",
51097=>X"00",
51098=>X"00",
51099=>X"00",
51100=>X"00",
51101=>X"00",
51102=>X"00",
51103=>X"00",
51104=>X"00",
51105=>X"00",
51106=>X"00",
51107=>X"00",
51108=>X"00",
51109=>X"00",
51110=>X"00",
51111=>X"00",
51112=>X"00",
51113=>X"00",
51114=>X"00",
51115=>X"00",
51116=>X"00",
51117=>X"00",
51118=>X"00",
51119=>X"00",
51120=>X"00",
51121=>X"00",
51122=>X"00",
51123=>X"00",
51124=>X"00",
51125=>X"00",
51126=>X"00",
51127=>X"00",
51128=>X"00",
51129=>X"00",
51130=>X"00",
51131=>X"00",
51132=>X"00",
51133=>X"00",
51134=>X"00",
51135=>X"00",
51136=>X"00",
51137=>X"00",
51138=>X"00",
51139=>X"00",
51140=>X"00",
51141=>X"00",
51142=>X"00",
51143=>X"00",
51144=>X"00",
51145=>X"00",
51146=>X"00",
51147=>X"00",
51148=>X"00",
51149=>X"00",
51150=>X"00",
51151=>X"00",
51152=>X"00",
51153=>X"00",
51154=>X"00",
51155=>X"00",
51156=>X"00",
51157=>X"00",
51158=>X"00",
51159=>X"00",
51160=>X"00",
51161=>X"00",
51162=>X"00",
51163=>X"00",
51164=>X"00",
51165=>X"00",
51166=>X"00",
51167=>X"00",
51168=>X"00",
51169=>X"00",
51170=>X"00",
51171=>X"00",
51172=>X"00",
51173=>X"00",
51174=>X"00",
51175=>X"00",
51176=>X"00",
51177=>X"00",
51178=>X"00",
51179=>X"00",
51180=>X"00",
51181=>X"00",
51182=>X"00",
51183=>X"00",
51184=>X"00",
51185=>X"00",
51186=>X"00",
51187=>X"00",
51188=>X"00",
51189=>X"00",
51190=>X"00",
51191=>X"00",
51192=>X"00",
51193=>X"00",
51194=>X"00",
51195=>X"00",
51196=>X"00",
51197=>X"00",
51198=>X"00",
51199=>X"00",
51200=>X"00",
51201=>X"00",
51202=>X"00",
51203=>X"00",
51204=>X"00",
51205=>X"00",
51206=>X"00",
51207=>X"00",
51208=>X"00",
51209=>X"00",
51210=>X"00",
51211=>X"00",
51212=>X"00",
51213=>X"00",
51214=>X"00",
51215=>X"00",
51216=>X"00",
51217=>X"00",
51218=>X"00",
51219=>X"00",
51220=>X"00",
51221=>X"00",
51222=>X"00",
51223=>X"00",
51224=>X"00",
51225=>X"00",
51226=>X"00",
51227=>X"00",
51228=>X"00",
51229=>X"00",
51230=>X"00",
51231=>X"00",
51232=>X"00",
51233=>X"00",
51234=>X"00",
51235=>X"00",
51236=>X"00",
51237=>X"00",
51238=>X"00",
51239=>X"00",
51240=>X"00",
51241=>X"00",
51242=>X"00",
51243=>X"00",
51244=>X"00",
51245=>X"00",
51246=>X"00",
51247=>X"00",
51248=>X"00",
51249=>X"00",
51250=>X"00",
51251=>X"00",
51252=>X"00",
51253=>X"00",
51254=>X"00",
51255=>X"00",
51256=>X"00",
51257=>X"00",
51258=>X"00",
51259=>X"00",
51260=>X"00",
51261=>X"00",
51262=>X"00",
51263=>X"00",
51264=>X"00",
51265=>X"00",
51266=>X"00",
51267=>X"00",
51268=>X"00",
51269=>X"00",
51270=>X"00",
51271=>X"00",
51272=>X"00",
51273=>X"00",
51274=>X"00",
51275=>X"00",
51276=>X"00",
51277=>X"00",
51278=>X"00",
51279=>X"00",
51280=>X"00",
51281=>X"00",
51282=>X"00",
51283=>X"00",
51284=>X"00",
51285=>X"00",
51286=>X"00",
51287=>X"00",
51288=>X"00",
51289=>X"00",
51290=>X"00",
51291=>X"00",
51292=>X"00",
51293=>X"00",
51294=>X"00",
51295=>X"00",
51296=>X"00",
51297=>X"00",
51298=>X"00",
51299=>X"00",
51300=>X"00",
51301=>X"00",
51302=>X"00",
51303=>X"00",
51304=>X"00",
51305=>X"00",
51306=>X"00",
51307=>X"00",
51308=>X"00",
51309=>X"00",
51310=>X"00",
51311=>X"00",
51312=>X"00",
51313=>X"00",
51314=>X"00",
51315=>X"00",
51316=>X"00",
51317=>X"00",
51318=>X"00",
51319=>X"00",
51320=>X"00",
51321=>X"00",
51322=>X"00",
51323=>X"00",
51324=>X"00",
51325=>X"00",
51326=>X"00",
51327=>X"00",
51328=>X"00",
51329=>X"00",
51330=>X"00",
51331=>X"00",
51332=>X"00",
51333=>X"00",
51334=>X"00",
51335=>X"00",
51336=>X"00",
51337=>X"00",
51338=>X"00",
51339=>X"00",
51340=>X"00",
51341=>X"00",
51342=>X"00",
51343=>X"00",
51344=>X"00",
51345=>X"00",
51346=>X"00",
51347=>X"00",
51348=>X"00",
51349=>X"00",
51350=>X"00",
51351=>X"00",
51352=>X"00",
51353=>X"00",
51354=>X"00",
51355=>X"00",
51356=>X"00",
51357=>X"00",
51358=>X"00",
51359=>X"00",
51360=>X"00",
51361=>X"00",
51362=>X"00",
51363=>X"00",
51364=>X"00",
51365=>X"00",
51366=>X"00",
51367=>X"00",
51368=>X"00",
51369=>X"00",
51370=>X"00",
51371=>X"00",
51372=>X"00",
51373=>X"00",
51374=>X"00",
51375=>X"00",
51376=>X"00",
51377=>X"00",
51378=>X"00",
51379=>X"00",
51380=>X"00",
51381=>X"00",
51382=>X"00",
51383=>X"00",
51384=>X"00",
51385=>X"00",
51386=>X"00",
51387=>X"00",
51388=>X"00",
51389=>X"00",
51390=>X"00",
51391=>X"00",
51392=>X"00",
51393=>X"00",
51394=>X"00",
51395=>X"00",
51396=>X"00",
51397=>X"00",
51398=>X"00",
51399=>X"00",
51400=>X"00",
51401=>X"00",
51402=>X"00",
51403=>X"00",
51404=>X"00",
51405=>X"00",
51406=>X"00",
51407=>X"00",
51408=>X"00",
51409=>X"00",
51410=>X"00",
51411=>X"00",
51412=>X"00",
51413=>X"00",
51414=>X"00",
51415=>X"00",
51416=>X"00",
51417=>X"00",
51418=>X"00",
51419=>X"00",
51420=>X"00",
51421=>X"00",
51422=>X"00",
51423=>X"00",
51424=>X"00",
51425=>X"00",
51426=>X"00",
51427=>X"00",
51428=>X"00",
51429=>X"00",
51430=>X"00",
51431=>X"00",
51432=>X"00",
51433=>X"00",
51434=>X"00",
51435=>X"00",
51436=>X"00",
51437=>X"00",
51438=>X"00",
51439=>X"00",
51440=>X"00",
51441=>X"00",
51442=>X"00",
51443=>X"00",
51444=>X"00",
51445=>X"00",
51446=>X"00",
51447=>X"00",
51448=>X"00",
51449=>X"00",
51450=>X"00",
51451=>X"00",
51452=>X"00",
51453=>X"00",
51454=>X"00",
51455=>X"00",
51456=>X"00",
51457=>X"00",
51458=>X"00",
51459=>X"00",
51460=>X"00",
51461=>X"00",
51462=>X"00",
51463=>X"00",
51464=>X"00",
51465=>X"00",
51466=>X"00",
51467=>X"00",
51468=>X"00",
51469=>X"00",
51470=>X"00",
51471=>X"00",
51472=>X"00",
51473=>X"00",
51474=>X"00",
51475=>X"00",
51476=>X"00",
51477=>X"00",
51478=>X"00",
51479=>X"00",
51480=>X"00",
51481=>X"00",
51482=>X"00",
51483=>X"00",
51484=>X"00",
51485=>X"00",
51486=>X"00",
51487=>X"00",
51488=>X"00",
51489=>X"00",
51490=>X"00",
51491=>X"00",
51492=>X"00",
51493=>X"00",
51494=>X"00",
51495=>X"00",
51496=>X"00",
51497=>X"00",
51498=>X"00",
51499=>X"00",
51500=>X"00",
51501=>X"00",
51502=>X"00",
51503=>X"00",
51504=>X"00",
51505=>X"00",
51506=>X"00",
51507=>X"00",
51508=>X"00",
51509=>X"00",
51510=>X"00",
51511=>X"00",
51512=>X"00",
51513=>X"00",
51514=>X"00",
51515=>X"00",
51516=>X"00",
51517=>X"00",
51518=>X"00",
51519=>X"00",
51520=>X"00",
51521=>X"00",
51522=>X"00",
51523=>X"00",
51524=>X"00",
51525=>X"00",
51526=>X"00",
51527=>X"00",
51528=>X"00",
51529=>X"00",
51530=>X"00",
51531=>X"00",
51532=>X"00",
51533=>X"00",
51534=>X"00",
51535=>X"00",
51536=>X"00",
51537=>X"00",
51538=>X"00",
51539=>X"00",
51540=>X"00",
51541=>X"00",
51542=>X"00",
51543=>X"00",
51544=>X"00",
51545=>X"00",
51546=>X"00",
51547=>X"00",
51548=>X"00",
51549=>X"00",
51550=>X"00",
51551=>X"00",
51552=>X"00",
51553=>X"00",
51554=>X"00",
51555=>X"00",
51556=>X"00",
51557=>X"00",
51558=>X"00",
51559=>X"00",
51560=>X"00",
51561=>X"00",
51562=>X"00",
51563=>X"00",
51564=>X"00",
51565=>X"00",
51566=>X"00",
51567=>X"00",
51568=>X"00",
51569=>X"00",
51570=>X"00",
51571=>X"00",
51572=>X"00",
51573=>X"00",
51574=>X"00",
51575=>X"00",
51576=>X"00",
51577=>X"00",
51578=>X"00",
51579=>X"00",
51580=>X"00",
51581=>X"00",
51582=>X"00",
51583=>X"00",
51584=>X"00",
51585=>X"00",
51586=>X"00",
51587=>X"00",
51588=>X"00",
51589=>X"00",
51590=>X"00",
51591=>X"00",
51592=>X"00",
51593=>X"00",
51594=>X"00",
51595=>X"00",
51596=>X"00",
51597=>X"00",
51598=>X"00",
51599=>X"00",
51600=>X"00",
51601=>X"00",
51602=>X"00",
51603=>X"00",
51604=>X"00",
51605=>X"00",
51606=>X"00",
51607=>X"00",
51608=>X"00",
51609=>X"00",
51610=>X"00",
51611=>X"00",
51612=>X"00",
51613=>X"00",
51614=>X"00",
51615=>X"00",
51616=>X"00",
51617=>X"00",
51618=>X"00",
51619=>X"00",
51620=>X"00",
51621=>X"00",
51622=>X"00",
51623=>X"00",
51624=>X"00",
51625=>X"00",
51626=>X"00",
51627=>X"00",
51628=>X"00",
51629=>X"00",
51630=>X"00",
51631=>X"00",
51632=>X"00",
51633=>X"00",
51634=>X"00",
51635=>X"00",
51636=>X"00",
51637=>X"00",
51638=>X"00",
51639=>X"00",
51640=>X"00",
51641=>X"00",
51642=>X"00",
51643=>X"00",
51644=>X"00",
51645=>X"00",
51646=>X"00",
51647=>X"00",
51648=>X"00",
51649=>X"00",
51650=>X"00",
51651=>X"00",
51652=>X"00",
51653=>X"00",
51654=>X"00",
51655=>X"00",
51656=>X"00",
51657=>X"00",
51658=>X"00",
51659=>X"00",
51660=>X"00",
51661=>X"00",
51662=>X"00",
51663=>X"00",
51664=>X"00",
51665=>X"00",
51666=>X"00",
51667=>X"00",
51668=>X"00",
51669=>X"00",
51670=>X"00",
51671=>X"00",
51672=>X"00",
51673=>X"00",
51674=>X"00",
51675=>X"00",
51676=>X"00",
51677=>X"00",
51678=>X"00",
51679=>X"00",
51680=>X"00",
51681=>X"00",
51682=>X"00",
51683=>X"00",
51684=>X"00",
51685=>X"00",
51686=>X"00",
51687=>X"00",
51688=>X"00",
51689=>X"00",
51690=>X"00",
51691=>X"00",
51692=>X"00",
51693=>X"00",
51694=>X"00",
51695=>X"00",
51696=>X"00",
51697=>X"00",
51698=>X"00",
51699=>X"00",
51700=>X"00",
51701=>X"00",
51702=>X"00",
51703=>X"00",
51704=>X"00",
51705=>X"00",
51706=>X"00",
51707=>X"00",
51708=>X"00",
51709=>X"00",
51710=>X"00",
51711=>X"00",
51712=>X"00",
51713=>X"00",
51714=>X"00",
51715=>X"00",
51716=>X"00",
51717=>X"00",
51718=>X"00",
51719=>X"00",
51720=>X"00",
51721=>X"00",
51722=>X"00",
51723=>X"00",
51724=>X"00",
51725=>X"00",
51726=>X"00",
51727=>X"00",
51728=>X"00",
51729=>X"00",
51730=>X"00",
51731=>X"00",
51732=>X"00",
51733=>X"00",
51734=>X"00",
51735=>X"00",
51736=>X"00",
51737=>X"00",
51738=>X"00",
51739=>X"00",
51740=>X"00",
51741=>X"00",
51742=>X"00",
51743=>X"00",
51744=>X"00",
51745=>X"00",
51746=>X"00",
51747=>X"00",
51748=>X"00",
51749=>X"00",
51750=>X"00",
51751=>X"00",
51752=>X"00",
51753=>X"00",
51754=>X"00",
51755=>X"00",
51756=>X"00",
51757=>X"00",
51758=>X"00",
51759=>X"00",
51760=>X"00",
51761=>X"00",
51762=>X"00",
51763=>X"00",
51764=>X"00",
51765=>X"00",
51766=>X"00",
51767=>X"00",
51768=>X"00",
51769=>X"00",
51770=>X"00",
51771=>X"00",
51772=>X"00",
51773=>X"00",
51774=>X"00",
51775=>X"00",
51776=>X"00",
51777=>X"00",
51778=>X"00",
51779=>X"00",
51780=>X"00",
51781=>X"00",
51782=>X"00",
51783=>X"00",
51784=>X"00",
51785=>X"00",
51786=>X"00",
51787=>X"00",
51788=>X"00",
51789=>X"00",
51790=>X"00",
51791=>X"00",
51792=>X"00",
51793=>X"00",
51794=>X"00",
51795=>X"00",
51796=>X"00",
51797=>X"00",
51798=>X"00",
51799=>X"00",
51800=>X"00",
51801=>X"00",
51802=>X"00",
51803=>X"00",
51804=>X"00",
51805=>X"00",
51806=>X"00",
51807=>X"00",
51808=>X"00",
51809=>X"00",
51810=>X"00",
51811=>X"00",
51812=>X"00",
51813=>X"00",
51814=>X"00",
51815=>X"00",
51816=>X"00",
51817=>X"00",
51818=>X"00",
51819=>X"00",
51820=>X"00",
51821=>X"00",
51822=>X"00",
51823=>X"00",
51824=>X"00",
51825=>X"00",
51826=>X"00",
51827=>X"00",
51828=>X"00",
51829=>X"00",
51830=>X"00",
51831=>X"00",
51832=>X"00",
51833=>X"00",
51834=>X"00",
51835=>X"00",
51836=>X"00",
51837=>X"00",
51838=>X"00",
51839=>X"00",
51840=>X"00",
51841=>X"00",
51842=>X"00",
51843=>X"00",
51844=>X"00",
51845=>X"00",
51846=>X"00",
51847=>X"00",
51848=>X"00",
51849=>X"00",
51850=>X"00",
51851=>X"00",
51852=>X"00",
51853=>X"00",
51854=>X"00",
51855=>X"00",
51856=>X"00",
51857=>X"00",
51858=>X"00",
51859=>X"00",
51860=>X"00",
51861=>X"00",
51862=>X"00",
51863=>X"00",
51864=>X"00",
51865=>X"00",
51866=>X"00",
51867=>X"00",
51868=>X"00",
51869=>X"00",
51870=>X"00",
51871=>X"00",
51872=>X"00",
51873=>X"00",
51874=>X"00",
51875=>X"00",
51876=>X"00",
51877=>X"00",
51878=>X"00",
51879=>X"00",
51880=>X"00",
51881=>X"00",
51882=>X"00",
51883=>X"00",
51884=>X"00",
51885=>X"00",
51886=>X"00",
51887=>X"00",
51888=>X"00",
51889=>X"00",
51890=>X"00",
51891=>X"00",
51892=>X"00",
51893=>X"00",
51894=>X"00",
51895=>X"00",
51896=>X"00",
51897=>X"00",
51898=>X"00",
51899=>X"00",
51900=>X"00",
51901=>X"00",
51902=>X"00",
51903=>X"00",
51904=>X"00",
51905=>X"00",
51906=>X"00",
51907=>X"00",
51908=>X"00",
51909=>X"00",
51910=>X"00",
51911=>X"00",
51912=>X"00",
51913=>X"00",
51914=>X"00",
51915=>X"00",
51916=>X"00",
51917=>X"00",
51918=>X"00",
51919=>X"00",
51920=>X"00",
51921=>X"00",
51922=>X"00",
51923=>X"00",
51924=>X"00",
51925=>X"00",
51926=>X"00",
51927=>X"00",
51928=>X"00",
51929=>X"00",
51930=>X"00",
51931=>X"00",
51932=>X"00",
51933=>X"00",
51934=>X"00",
51935=>X"00",
51936=>X"00",
51937=>X"00",
51938=>X"00",
51939=>X"00",
51940=>X"00",
51941=>X"00",
51942=>X"00",
51943=>X"00",
51944=>X"00",
51945=>X"00",
51946=>X"00",
51947=>X"00",
51948=>X"00",
51949=>X"00",
51950=>X"00",
51951=>X"00",
51952=>X"00",
51953=>X"00",
51954=>X"00",
51955=>X"00",
51956=>X"00",
51957=>X"00",
51958=>X"00",
51959=>X"00",
51960=>X"00",
51961=>X"00",
51962=>X"00",
51963=>X"00",
51964=>X"00",
51965=>X"00",
51966=>X"00",
51967=>X"00",
51968=>X"00",
51969=>X"00",
51970=>X"00",
51971=>X"00",
51972=>X"00",
51973=>X"00",
51974=>X"00",
51975=>X"00",
51976=>X"00",
51977=>X"00",
51978=>X"00",
51979=>X"00",
51980=>X"00",
51981=>X"00",
51982=>X"00",
51983=>X"00",
51984=>X"00",
51985=>X"00",
51986=>X"00",
51987=>X"00",
51988=>X"00",
51989=>X"00",
51990=>X"00",
51991=>X"00",
51992=>X"00",
51993=>X"00",
51994=>X"00",
51995=>X"00",
51996=>X"00",
51997=>X"00",
51998=>X"00",
51999=>X"00",
52000=>X"00",
52001=>X"00",
52002=>X"00",
52003=>X"00",
52004=>X"00",
52005=>X"00",
52006=>X"00",
52007=>X"00",
52008=>X"00",
52009=>X"00",
52010=>X"00",
52011=>X"00",
52012=>X"00",
52013=>X"00",
52014=>X"00",
52015=>X"00",
52016=>X"00",
52017=>X"00",
52018=>X"00",
52019=>X"00",
52020=>X"00",
52021=>X"00",
52022=>X"00",
52023=>X"00",
52024=>X"00",
52025=>X"00",
52026=>X"00",
52027=>X"00",
52028=>X"00",
52029=>X"00",
52030=>X"00",
52031=>X"00",
52032=>X"00",
52033=>X"00",
52034=>X"00",
52035=>X"00",
52036=>X"00",
52037=>X"00",
52038=>X"00",
52039=>X"00",
52040=>X"00",
52041=>X"00",
52042=>X"00",
52043=>X"00",
52044=>X"00",
52045=>X"00",
52046=>X"00",
52047=>X"00",
52048=>X"00",
52049=>X"00",
52050=>X"00",
52051=>X"00",
52052=>X"00",
52053=>X"00",
52054=>X"00",
52055=>X"00",
52056=>X"00",
52057=>X"00",
52058=>X"00",
52059=>X"00",
52060=>X"00",
52061=>X"00",
52062=>X"00",
52063=>X"00",
52064=>X"00",
52065=>X"00",
52066=>X"00",
52067=>X"00",
52068=>X"00",
52069=>X"00",
52070=>X"00",
52071=>X"00",
52072=>X"00",
52073=>X"00",
52074=>X"00",
52075=>X"00",
52076=>X"00",
52077=>X"00",
52078=>X"00",
52079=>X"00",
52080=>X"00",
52081=>X"00",
52082=>X"00",
52083=>X"00",
52084=>X"00",
52085=>X"00",
52086=>X"00",
52087=>X"00",
52088=>X"00",
52089=>X"00",
52090=>X"00",
52091=>X"00",
52092=>X"00",
52093=>X"00",
52094=>X"00",
52095=>X"00",
52096=>X"00",
52097=>X"00",
52098=>X"00",
52099=>X"00",
52100=>X"00",
52101=>X"00",
52102=>X"00",
52103=>X"00",
52104=>X"00",
52105=>X"00",
52106=>X"00",
52107=>X"00",
52108=>X"00",
52109=>X"00",
52110=>X"00",
52111=>X"00",
52112=>X"00",
52113=>X"00",
52114=>X"00",
52115=>X"00",
52116=>X"00",
52117=>X"00",
52118=>X"00",
52119=>X"00",
52120=>X"00",
52121=>X"00",
52122=>X"00",
52123=>X"00",
52124=>X"00",
52125=>X"00",
52126=>X"00",
52127=>X"00",
52128=>X"00",
52129=>X"00",
52130=>X"00",
52131=>X"00",
52132=>X"00",
52133=>X"00",
52134=>X"00",
52135=>X"00",
52136=>X"00",
52137=>X"00",
52138=>X"00",
52139=>X"00",
52140=>X"00",
52141=>X"00",
52142=>X"00",
52143=>X"00",
52144=>X"00",
52145=>X"00",
52146=>X"00",
52147=>X"00",
52148=>X"00",
52149=>X"00",
52150=>X"00",
52151=>X"00",
52152=>X"00",
52153=>X"00",
52154=>X"00",
52155=>X"00",
52156=>X"00",
52157=>X"00",
52158=>X"00",
52159=>X"00",
52160=>X"00",
52161=>X"00",
52162=>X"00",
52163=>X"00",
52164=>X"00",
52165=>X"00",
52166=>X"00",
52167=>X"00",
52168=>X"00",
52169=>X"00",
52170=>X"00",
52171=>X"00",
52172=>X"00",
52173=>X"00",
52174=>X"00",
52175=>X"00",
52176=>X"00",
52177=>X"00",
52178=>X"00",
52179=>X"00",
52180=>X"00",
52181=>X"00",
52182=>X"00",
52183=>X"00",
52184=>X"00",
52185=>X"00",
52186=>X"00",
52187=>X"00",
52188=>X"00",
52189=>X"00",
52190=>X"00",
52191=>X"00",
52192=>X"00",
52193=>X"00",
52194=>X"00",
52195=>X"00",
52196=>X"00",
52197=>X"00",
52198=>X"00",
52199=>X"00",
52200=>X"00",
52201=>X"00",
52202=>X"00",
52203=>X"00",
52204=>X"00",
52205=>X"00",
52206=>X"00",
52207=>X"00",
52208=>X"00",
52209=>X"00",
52210=>X"00",
52211=>X"00",
52212=>X"00",
52213=>X"00",
52214=>X"00",
52215=>X"00",
52216=>X"00",
52217=>X"00",
52218=>X"00",
52219=>X"00",
52220=>X"00",
52221=>X"00",
52222=>X"00",
52223=>X"00",
52224=>X"00",
52225=>X"00",
52226=>X"00",
52227=>X"00",
52228=>X"00",
52229=>X"00",
52230=>X"00",
52231=>X"00",
52232=>X"00",
52233=>X"00",
52234=>X"00",
52235=>X"00",
52236=>X"00",
52237=>X"00",
52238=>X"00",
52239=>X"00",
52240=>X"00",
52241=>X"00",
52242=>X"00",
52243=>X"00",
52244=>X"00",
52245=>X"00",
52246=>X"00",
52247=>X"00",
52248=>X"00",
52249=>X"00",
52250=>X"00",
52251=>X"00",
52252=>X"00",
52253=>X"00",
52254=>X"00",
52255=>X"00",
52256=>X"00",
52257=>X"00",
52258=>X"00",
52259=>X"00",
52260=>X"00",
52261=>X"00",
52262=>X"00",
52263=>X"00",
52264=>X"00",
52265=>X"00",
52266=>X"00",
52267=>X"00",
52268=>X"00",
52269=>X"00",
52270=>X"00",
52271=>X"00",
52272=>X"00",
52273=>X"00",
52274=>X"00",
52275=>X"00",
52276=>X"00",
52277=>X"00",
52278=>X"00",
52279=>X"00",
52280=>X"00",
52281=>X"00",
52282=>X"00",
52283=>X"00",
52284=>X"00",
52285=>X"00",
52286=>X"00",
52287=>X"00",
52288=>X"00",
52289=>X"00",
52290=>X"00",
52291=>X"00",
52292=>X"00",
52293=>X"00",
52294=>X"00",
52295=>X"00",
52296=>X"00",
52297=>X"00",
52298=>X"00",
52299=>X"00",
52300=>X"00",
52301=>X"00",
52302=>X"00",
52303=>X"00",
52304=>X"00",
52305=>X"00",
52306=>X"00",
52307=>X"00",
52308=>X"00",
52309=>X"00",
52310=>X"00",
52311=>X"00",
52312=>X"00",
52313=>X"00",
52314=>X"00",
52315=>X"00",
52316=>X"00",
52317=>X"00",
52318=>X"00",
52319=>X"00",
52320=>X"00",
52321=>X"00",
52322=>X"00",
52323=>X"00",
52324=>X"00",
52325=>X"00",
52326=>X"00",
52327=>X"00",
52328=>X"00",
52329=>X"00",
52330=>X"00",
52331=>X"00",
52332=>X"00",
52333=>X"00",
52334=>X"00",
52335=>X"00",
52336=>X"00",
52337=>X"00",
52338=>X"00",
52339=>X"00",
52340=>X"00",
52341=>X"00",
52342=>X"00",
52343=>X"00",
52344=>X"00",
52345=>X"00",
52346=>X"00",
52347=>X"00",
52348=>X"00",
52349=>X"00",
52350=>X"00",
52351=>X"00",
52352=>X"00",
52353=>X"00",
52354=>X"00",
52355=>X"00",
52356=>X"00",
52357=>X"00",
52358=>X"00",
52359=>X"00",
52360=>X"00",
52361=>X"00",
52362=>X"00",
52363=>X"00",
52364=>X"00",
52365=>X"00",
52366=>X"00",
52367=>X"00",
52368=>X"00",
52369=>X"00",
52370=>X"00",
52371=>X"00",
52372=>X"00",
52373=>X"00",
52374=>X"00",
52375=>X"00",
52376=>X"00",
52377=>X"00",
52378=>X"00",
52379=>X"00",
52380=>X"00",
52381=>X"00",
52382=>X"00",
52383=>X"00",
52384=>X"00",
52385=>X"00",
52386=>X"00",
52387=>X"00",
52388=>X"00",
52389=>X"00",
52390=>X"00",
52391=>X"00",
52392=>X"00",
52393=>X"00",
52394=>X"00",
52395=>X"00",
52396=>X"00",
52397=>X"00",
52398=>X"00",
52399=>X"00",
52400=>X"00",
52401=>X"00",
52402=>X"00",
52403=>X"00",
52404=>X"00",
52405=>X"00",
52406=>X"00",
52407=>X"00",
52408=>X"00",
52409=>X"00",
52410=>X"00",
52411=>X"00",
52412=>X"00",
52413=>X"00",
52414=>X"00",
52415=>X"00",
52416=>X"00",
52417=>X"00",
52418=>X"00",
52419=>X"00",
52420=>X"00",
52421=>X"00",
52422=>X"00",
52423=>X"00",
52424=>X"00",
52425=>X"00",
52426=>X"00",
52427=>X"00",
52428=>X"00",
52429=>X"00",
52430=>X"00",
52431=>X"00",
52432=>X"00",
52433=>X"00",
52434=>X"00",
52435=>X"00",
52436=>X"00",
52437=>X"00",
52438=>X"00",
52439=>X"00",
52440=>X"00",
52441=>X"00",
52442=>X"00",
52443=>X"00",
52444=>X"00",
52445=>X"00",
52446=>X"00",
52447=>X"00",
52448=>X"00",
52449=>X"00",
52450=>X"00",
52451=>X"00",
52452=>X"00",
52453=>X"00",
52454=>X"00",
52455=>X"00",
52456=>X"00",
52457=>X"00",
52458=>X"00",
52459=>X"00",
52460=>X"00",
52461=>X"00",
52462=>X"00",
52463=>X"00",
52464=>X"00",
52465=>X"00",
52466=>X"00",
52467=>X"00",
52468=>X"00",
52469=>X"00",
52470=>X"00",
52471=>X"00",
52472=>X"00",
52473=>X"00",
52474=>X"00",
52475=>X"00",
52476=>X"00",
52477=>X"00",
52478=>X"00",
52479=>X"00",
52480=>X"00",
52481=>X"00",
52482=>X"00",
52483=>X"00",
52484=>X"00",
52485=>X"00",
52486=>X"00",
52487=>X"00",
52488=>X"00",
52489=>X"00",
52490=>X"00",
52491=>X"00",
52492=>X"00",
52493=>X"00",
52494=>X"00",
52495=>X"00",
52496=>X"00",
52497=>X"00",
52498=>X"00",
52499=>X"00",
52500=>X"00",
52501=>X"00",
52502=>X"00",
52503=>X"00",
52504=>X"00",
52505=>X"00",
52506=>X"00",
52507=>X"00",
52508=>X"00",
52509=>X"00",
52510=>X"00",
52511=>X"00",
52512=>X"00",
52513=>X"00",
52514=>X"00",
52515=>X"00",
52516=>X"00",
52517=>X"00",
52518=>X"00",
52519=>X"00",
52520=>X"00",
52521=>X"00",
52522=>X"00",
52523=>X"00",
52524=>X"00",
52525=>X"00",
52526=>X"00",
52527=>X"00",
52528=>X"00",
52529=>X"00",
52530=>X"00",
52531=>X"00",
52532=>X"00",
52533=>X"00",
52534=>X"00",
52535=>X"00",
52536=>X"00",
52537=>X"00",
52538=>X"00",
52539=>X"00",
52540=>X"00",
52541=>X"00",
52542=>X"00",
52543=>X"00",
52544=>X"00",
52545=>X"00",
52546=>X"00",
52547=>X"00",
52548=>X"00",
52549=>X"00",
52550=>X"00",
52551=>X"00",
52552=>X"00",
52553=>X"00",
52554=>X"00",
52555=>X"00",
52556=>X"00",
52557=>X"00",
52558=>X"00",
52559=>X"00",
52560=>X"00",
52561=>X"00",
52562=>X"00",
52563=>X"00",
52564=>X"00",
52565=>X"00",
52566=>X"00",
52567=>X"00",
52568=>X"00",
52569=>X"00",
52570=>X"00",
52571=>X"00",
52572=>X"00",
52573=>X"00",
52574=>X"00",
52575=>X"00",
52576=>X"00",
52577=>X"00",
52578=>X"00",
52579=>X"00",
52580=>X"00",
52581=>X"00",
52582=>X"00",
52583=>X"00",
52584=>X"00",
52585=>X"00",
52586=>X"00",
52587=>X"00",
52588=>X"00",
52589=>X"00",
52590=>X"00",
52591=>X"00",
52592=>X"00",
52593=>X"00",
52594=>X"00",
52595=>X"00",
52596=>X"00",
52597=>X"00",
52598=>X"00",
52599=>X"00",
52600=>X"00",
52601=>X"00",
52602=>X"00",
52603=>X"00",
52604=>X"00",
52605=>X"00",
52606=>X"00",
52607=>X"00",
52608=>X"00",
52609=>X"00",
52610=>X"00",
52611=>X"00",
52612=>X"00",
52613=>X"00",
52614=>X"00",
52615=>X"00",
52616=>X"00",
52617=>X"00",
52618=>X"00",
52619=>X"00",
52620=>X"00",
52621=>X"00",
52622=>X"00",
52623=>X"00",
52624=>X"00",
52625=>X"00",
52626=>X"00",
52627=>X"00",
52628=>X"00",
52629=>X"00",
52630=>X"00",
52631=>X"00",
52632=>X"00",
52633=>X"00",
52634=>X"00",
52635=>X"00",
52636=>X"00",
52637=>X"00",
52638=>X"00",
52639=>X"00",
52640=>X"00",
52641=>X"00",
52642=>X"00",
52643=>X"00",
52644=>X"00",
52645=>X"00",
52646=>X"00",
52647=>X"00",
52648=>X"00",
52649=>X"00",
52650=>X"00",
52651=>X"00",
52652=>X"00",
52653=>X"00",
52654=>X"00",
52655=>X"00",
52656=>X"00",
52657=>X"00",
52658=>X"00",
52659=>X"00",
52660=>X"00",
52661=>X"00",
52662=>X"00",
52663=>X"00",
52664=>X"00",
52665=>X"00",
52666=>X"00",
52667=>X"00",
52668=>X"00",
52669=>X"00",
52670=>X"00",
52671=>X"00",
52672=>X"00",
52673=>X"00",
52674=>X"00",
52675=>X"00",
52676=>X"00",
52677=>X"00",
52678=>X"00",
52679=>X"00",
52680=>X"00",
52681=>X"00",
52682=>X"00",
52683=>X"00",
52684=>X"00",
52685=>X"00",
52686=>X"00",
52687=>X"00",
52688=>X"00",
52689=>X"00",
52690=>X"00",
52691=>X"00",
52692=>X"00",
52693=>X"00",
52694=>X"00",
52695=>X"00",
52696=>X"00",
52697=>X"00",
52698=>X"00",
52699=>X"00",
52700=>X"00",
52701=>X"00",
52702=>X"00",
52703=>X"00",
52704=>X"00",
52705=>X"00",
52706=>X"00",
52707=>X"00",
52708=>X"00",
52709=>X"00",
52710=>X"00",
52711=>X"00",
52712=>X"00",
52713=>X"00",
52714=>X"00",
52715=>X"00",
52716=>X"00",
52717=>X"00",
52718=>X"00",
52719=>X"00",
52720=>X"00",
52721=>X"00",
52722=>X"00",
52723=>X"00",
52724=>X"00",
52725=>X"00",
52726=>X"00",
52727=>X"00",
52728=>X"00",
52729=>X"00",
52730=>X"00",
52731=>X"00",
52732=>X"00",
52733=>X"00",
52734=>X"00",
52735=>X"00",
52736=>X"00",
52737=>X"00",
52738=>X"00",
52739=>X"00",
52740=>X"00",
52741=>X"00",
52742=>X"00",
52743=>X"00",
52744=>X"00",
52745=>X"00",
52746=>X"00",
52747=>X"00",
52748=>X"00",
52749=>X"00",
52750=>X"00",
52751=>X"00",
52752=>X"00",
52753=>X"00",
52754=>X"00",
52755=>X"00",
52756=>X"00",
52757=>X"00",
52758=>X"00",
52759=>X"00",
52760=>X"00",
52761=>X"00",
52762=>X"00",
52763=>X"00",
52764=>X"00",
52765=>X"00",
52766=>X"00",
52767=>X"00",
52768=>X"00",
52769=>X"00",
52770=>X"00",
52771=>X"00",
52772=>X"00",
52773=>X"00",
52774=>X"00",
52775=>X"00",
52776=>X"00",
52777=>X"00",
52778=>X"00",
52779=>X"00",
52780=>X"00",
52781=>X"00",
52782=>X"00",
52783=>X"00",
52784=>X"00",
52785=>X"00",
52786=>X"00",
52787=>X"00",
52788=>X"00",
52789=>X"00",
52790=>X"00",
52791=>X"00",
52792=>X"00",
52793=>X"00",
52794=>X"00",
52795=>X"00",
52796=>X"00",
52797=>X"00",
52798=>X"00",
52799=>X"00",
52800=>X"00",
52801=>X"00",
52802=>X"00",
52803=>X"00",
52804=>X"00",
52805=>X"00",
52806=>X"00",
52807=>X"00",
52808=>X"00",
52809=>X"00",
52810=>X"00",
52811=>X"00",
52812=>X"00",
52813=>X"00",
52814=>X"00",
52815=>X"00",
52816=>X"00",
52817=>X"00",
52818=>X"00",
52819=>X"00",
52820=>X"00",
52821=>X"00",
52822=>X"00",
52823=>X"00",
52824=>X"00",
52825=>X"00",
52826=>X"00",
52827=>X"00",
52828=>X"00",
52829=>X"00",
52830=>X"00",
52831=>X"00",
52832=>X"00",
52833=>X"00",
52834=>X"00",
52835=>X"00",
52836=>X"00",
52837=>X"00",
52838=>X"00",
52839=>X"00",
52840=>X"00",
52841=>X"00",
52842=>X"00",
52843=>X"00",
52844=>X"00",
52845=>X"00",
52846=>X"00",
52847=>X"00",
52848=>X"00",
52849=>X"00",
52850=>X"00",
52851=>X"00",
52852=>X"00",
52853=>X"00",
52854=>X"00",
52855=>X"00",
52856=>X"00",
52857=>X"00",
52858=>X"00",
52859=>X"00",
52860=>X"00",
52861=>X"00",
52862=>X"00",
52863=>X"00",
52864=>X"00",
52865=>X"00",
52866=>X"00",
52867=>X"00",
52868=>X"00",
52869=>X"00",
52870=>X"00",
52871=>X"00",
52872=>X"00",
52873=>X"00",
52874=>X"00",
52875=>X"00",
52876=>X"00",
52877=>X"00",
52878=>X"00",
52879=>X"00",
52880=>X"00",
52881=>X"00",
52882=>X"00",
52883=>X"00",
52884=>X"00",
52885=>X"00",
52886=>X"00",
52887=>X"00",
52888=>X"00",
52889=>X"00",
52890=>X"00",
52891=>X"00",
52892=>X"00",
52893=>X"00",
52894=>X"00",
52895=>X"00",
52896=>X"00",
52897=>X"00",
52898=>X"00",
52899=>X"00",
52900=>X"00",
52901=>X"00",
52902=>X"00",
52903=>X"00",
52904=>X"00",
52905=>X"00",
52906=>X"00",
52907=>X"00",
52908=>X"00",
52909=>X"00",
52910=>X"00",
52911=>X"00",
52912=>X"00",
52913=>X"00",
52914=>X"00",
52915=>X"00",
52916=>X"00",
52917=>X"00",
52918=>X"00",
52919=>X"00",
52920=>X"00",
52921=>X"00",
52922=>X"00",
52923=>X"00",
52924=>X"00",
52925=>X"00",
52926=>X"00",
52927=>X"00",
52928=>X"00",
52929=>X"00",
52930=>X"00",
52931=>X"00",
52932=>X"00",
52933=>X"00",
52934=>X"00",
52935=>X"00",
52936=>X"00",
52937=>X"00",
52938=>X"00",
52939=>X"00",
52940=>X"00",
52941=>X"00",
52942=>X"00",
52943=>X"00",
52944=>X"00",
52945=>X"00",
52946=>X"00",
52947=>X"00",
52948=>X"00",
52949=>X"00",
52950=>X"00",
52951=>X"00",
52952=>X"00",
52953=>X"00",
52954=>X"00",
52955=>X"00",
52956=>X"00",
52957=>X"00",
52958=>X"00",
52959=>X"00",
52960=>X"00",
52961=>X"00",
52962=>X"00",
52963=>X"00",
52964=>X"00",
52965=>X"00",
52966=>X"00",
52967=>X"00",
52968=>X"00",
52969=>X"00",
52970=>X"00",
52971=>X"00",
52972=>X"00",
52973=>X"00",
52974=>X"00",
52975=>X"00",
52976=>X"00",
52977=>X"00",
52978=>X"00",
52979=>X"00",
52980=>X"00",
52981=>X"00",
52982=>X"00",
52983=>X"00",
52984=>X"00",
52985=>X"00",
52986=>X"00",
52987=>X"00",
52988=>X"00",
52989=>X"00",
52990=>X"00",
52991=>X"00",
52992=>X"00",
52993=>X"00",
52994=>X"00",
52995=>X"00",
52996=>X"00",
52997=>X"00",
52998=>X"00",
52999=>X"00",
53000=>X"00",
53001=>X"00",
53002=>X"00",
53003=>X"00",
53004=>X"00",
53005=>X"00",
53006=>X"00",
53007=>X"00",
53008=>X"00",
53009=>X"00",
53010=>X"00",
53011=>X"00",
53012=>X"00",
53013=>X"00",
53014=>X"00",
53015=>X"00",
53016=>X"00",
53017=>X"00",
53018=>X"00",
53019=>X"00",
53020=>X"00",
53021=>X"00",
53022=>X"00",
53023=>X"00",
53024=>X"00",
53025=>X"00",
53026=>X"00",
53027=>X"00",
53028=>X"00",
53029=>X"00",
53030=>X"00",
53031=>X"00",
53032=>X"00",
53033=>X"00",
53034=>X"00",
53035=>X"00",
53036=>X"00",
53037=>X"00",
53038=>X"00",
53039=>X"00",
53040=>X"00",
53041=>X"00",
53042=>X"00",
53043=>X"00",
53044=>X"00",
53045=>X"00",
53046=>X"00",
53047=>X"00",
53048=>X"00",
53049=>X"00",
53050=>X"00",
53051=>X"00",
53052=>X"00",
53053=>X"00",
53054=>X"00",
53055=>X"00",
53056=>X"00",
53057=>X"00",
53058=>X"00",
53059=>X"00",
53060=>X"00",
53061=>X"00",
53062=>X"00",
53063=>X"00",
53064=>X"00",
53065=>X"00",
53066=>X"00",
53067=>X"00",
53068=>X"00",
53069=>X"00",
53070=>X"00",
53071=>X"00",
53072=>X"00",
53073=>X"00",
53074=>X"00",
53075=>X"00",
53076=>X"00",
53077=>X"00",
53078=>X"00",
53079=>X"00",
53080=>X"00",
53081=>X"00",
53082=>X"00",
53083=>X"00",
53084=>X"00",
53085=>X"00",
53086=>X"00",
53087=>X"00",
53088=>X"00",
53089=>X"00",
53090=>X"00",
53091=>X"00",
53092=>X"00",
53093=>X"00",
53094=>X"00",
53095=>X"00",
53096=>X"00",
53097=>X"00",
53098=>X"00",
53099=>X"00",
53100=>X"00",
53101=>X"00",
53102=>X"00",
53103=>X"00",
53104=>X"00",
53105=>X"00",
53106=>X"00",
53107=>X"00",
53108=>X"00",
53109=>X"00",
53110=>X"00",
53111=>X"00",
53112=>X"00",
53113=>X"00",
53114=>X"00",
53115=>X"00",
53116=>X"00",
53117=>X"00",
53118=>X"00",
53119=>X"00",
53120=>X"00",
53121=>X"00",
53122=>X"00",
53123=>X"00",
53124=>X"00",
53125=>X"00",
53126=>X"00",
53127=>X"00",
53128=>X"00",
53129=>X"00",
53130=>X"00",
53131=>X"00",
53132=>X"00",
53133=>X"00",
53134=>X"00",
53135=>X"00",
53136=>X"00",
53137=>X"00",
53138=>X"00",
53139=>X"00",
53140=>X"00",
53141=>X"00",
53142=>X"00",
53143=>X"00",
53144=>X"00",
53145=>X"00",
53146=>X"00",
53147=>X"00",
53148=>X"00",
53149=>X"00",
53150=>X"00",
53151=>X"00",
53152=>X"00",
53153=>X"00",
53154=>X"00",
53155=>X"00",
53156=>X"00",
53157=>X"00",
53158=>X"00",
53159=>X"00",
53160=>X"00",
53161=>X"00",
53162=>X"00",
53163=>X"00",
53164=>X"00",
53165=>X"00",
53166=>X"00",
53167=>X"00",
53168=>X"00",
53169=>X"00",
53170=>X"00",
53171=>X"00",
53172=>X"00",
53173=>X"00",
53174=>X"00",
53175=>X"00",
53176=>X"00",
53177=>X"00",
53178=>X"00",
53179=>X"00",
53180=>X"00",
53181=>X"00",
53182=>X"00",
53183=>X"00",
53184=>X"00",
53185=>X"00",
53186=>X"00",
53187=>X"00",
53188=>X"00",
53189=>X"00",
53190=>X"00",
53191=>X"00",
53192=>X"00",
53193=>X"00",
53194=>X"00",
53195=>X"00",
53196=>X"00",
53197=>X"00",
53198=>X"00",
53199=>X"00",
53200=>X"00",
53201=>X"00",
53202=>X"00",
53203=>X"00",
53204=>X"00",
53205=>X"00",
53206=>X"00",
53207=>X"00",
53208=>X"00",
53209=>X"00",
53210=>X"00",
53211=>X"00",
53212=>X"00",
53213=>X"00",
53214=>X"00",
53215=>X"00",
53216=>X"00",
53217=>X"00",
53218=>X"00",
53219=>X"00",
53220=>X"00",
53221=>X"00",
53222=>X"00",
53223=>X"00",
53224=>X"00",
53225=>X"00",
53226=>X"00",
53227=>X"00",
53228=>X"00",
53229=>X"00",
53230=>X"00",
53231=>X"00",
53232=>X"00",
53233=>X"00",
53234=>X"00",
53235=>X"00",
53236=>X"00",
53237=>X"00",
53238=>X"00",
53239=>X"00",
53240=>X"00",
53241=>X"00",
53242=>X"00",
53243=>X"00",
53244=>X"00",
53245=>X"00",
53246=>X"00",
53247=>X"00",
53248=>X"00",
53249=>X"00",
53250=>X"00",
53251=>X"00",
53252=>X"00",
53253=>X"00",
53254=>X"00",
53255=>X"00",
53256=>X"00",
53257=>X"00",
53258=>X"00",
53259=>X"00",
53260=>X"00",
53261=>X"00",
53262=>X"00",
53263=>X"00",
53264=>X"00",
53265=>X"00",
53266=>X"00",
53267=>X"00",
53268=>X"00",
53269=>X"00",
53270=>X"00",
53271=>X"00",
53272=>X"00",
53273=>X"00",
53274=>X"00",
53275=>X"00",
53276=>X"00",
53277=>X"00",
53278=>X"00",
53279=>X"00",
53280=>X"00",
53281=>X"00",
53282=>X"00",
53283=>X"00",
53284=>X"00",
53285=>X"00",
53286=>X"00",
53287=>X"00",
53288=>X"00",
53289=>X"00",
53290=>X"00",
53291=>X"00",
53292=>X"00",
53293=>X"00",
53294=>X"00",
53295=>X"00",
53296=>X"00",
53297=>X"00",
53298=>X"00",
53299=>X"00",
53300=>X"00",
53301=>X"00",
53302=>X"00",
53303=>X"00",
53304=>X"00",
53305=>X"00",
53306=>X"00",
53307=>X"00",
53308=>X"00",
53309=>X"00",
53310=>X"00",
53311=>X"00",
53312=>X"00",
53313=>X"00",
53314=>X"00",
53315=>X"00",
53316=>X"00",
53317=>X"00",
53318=>X"00",
53319=>X"00",
53320=>X"00",
53321=>X"00",
53322=>X"00",
53323=>X"00",
53324=>X"00",
53325=>X"00",
53326=>X"00",
53327=>X"00",
53328=>X"00",
53329=>X"00",
53330=>X"00",
53331=>X"00",
53332=>X"00",
53333=>X"00",
53334=>X"00",
53335=>X"00",
53336=>X"00",
53337=>X"00",
53338=>X"00",
53339=>X"00",
53340=>X"00",
53341=>X"00",
53342=>X"00",
53343=>X"00",
53344=>X"00",
53345=>X"00",
53346=>X"00",
53347=>X"00",
53348=>X"00",
53349=>X"00",
53350=>X"00",
53351=>X"00",
53352=>X"00",
53353=>X"00",
53354=>X"00",
53355=>X"00",
53356=>X"00",
53357=>X"00",
53358=>X"00",
53359=>X"00",
53360=>X"00",
53361=>X"00",
53362=>X"00",
53363=>X"00",
53364=>X"00",
53365=>X"00",
53366=>X"00",
53367=>X"00",
53368=>X"00",
53369=>X"00",
53370=>X"00",
53371=>X"00",
53372=>X"00",
53373=>X"00",
53374=>X"00",
53375=>X"00",
53376=>X"00",
53377=>X"00",
53378=>X"00",
53379=>X"00",
53380=>X"00",
53381=>X"00",
53382=>X"00",
53383=>X"00",
53384=>X"00",
53385=>X"00",
53386=>X"00",
53387=>X"00",
53388=>X"00",
53389=>X"00",
53390=>X"00",
53391=>X"00",
53392=>X"00",
53393=>X"00",
53394=>X"00",
53395=>X"00",
53396=>X"00",
53397=>X"00",
53398=>X"00",
53399=>X"00",
53400=>X"00",
53401=>X"00",
53402=>X"00",
53403=>X"00",
53404=>X"00",
53405=>X"00",
53406=>X"00",
53407=>X"00",
53408=>X"00",
53409=>X"00",
53410=>X"00",
53411=>X"00",
53412=>X"00",
53413=>X"00",
53414=>X"00",
53415=>X"00",
53416=>X"00",
53417=>X"00",
53418=>X"00",
53419=>X"00",
53420=>X"00",
53421=>X"00",
53422=>X"00",
53423=>X"00",
53424=>X"00",
53425=>X"00",
53426=>X"00",
53427=>X"00",
53428=>X"00",
53429=>X"00",
53430=>X"00",
53431=>X"00",
53432=>X"00",
53433=>X"00",
53434=>X"00",
53435=>X"00",
53436=>X"00",
53437=>X"00",
53438=>X"00",
53439=>X"00",
53440=>X"00",
53441=>X"00",
53442=>X"00",
53443=>X"00",
53444=>X"00",
53445=>X"00",
53446=>X"00",
53447=>X"00",
53448=>X"00",
53449=>X"00",
53450=>X"00",
53451=>X"00",
53452=>X"00",
53453=>X"00",
53454=>X"00",
53455=>X"00",
53456=>X"00",
53457=>X"00",
53458=>X"00",
53459=>X"00",
53460=>X"00",
53461=>X"00",
53462=>X"00",
53463=>X"00",
53464=>X"00",
53465=>X"00",
53466=>X"00",
53467=>X"00",
53468=>X"00",
53469=>X"00",
53470=>X"00",
53471=>X"00",
53472=>X"00",
53473=>X"00",
53474=>X"00",
53475=>X"00",
53476=>X"00",
53477=>X"00",
53478=>X"00",
53479=>X"00",
53480=>X"00",
53481=>X"00",
53482=>X"00",
53483=>X"00",
53484=>X"00",
53485=>X"00",
53486=>X"00",
53487=>X"00",
53488=>X"00",
53489=>X"00",
53490=>X"00",
53491=>X"00",
53492=>X"00",
53493=>X"00",
53494=>X"00",
53495=>X"00",
53496=>X"00",
53497=>X"00",
53498=>X"00",
53499=>X"00",
53500=>X"00",
53501=>X"00",
53502=>X"00",
53503=>X"00",
53504=>X"00",
53505=>X"00",
53506=>X"00",
53507=>X"00",
53508=>X"00",
53509=>X"00",
53510=>X"00",
53511=>X"00",
53512=>X"00",
53513=>X"00",
53514=>X"00",
53515=>X"00",
53516=>X"00",
53517=>X"00",
53518=>X"00",
53519=>X"00",
53520=>X"00",
53521=>X"00",
53522=>X"00",
53523=>X"00",
53524=>X"00",
53525=>X"00",
53526=>X"00",
53527=>X"00",
53528=>X"00",
53529=>X"00",
53530=>X"00",
53531=>X"00",
53532=>X"00",
53533=>X"00",
53534=>X"00",
53535=>X"00",
53536=>X"00",
53537=>X"00",
53538=>X"00",
53539=>X"00",
53540=>X"00",
53541=>X"00",
53542=>X"00",
53543=>X"00",
53544=>X"00",
53545=>X"00",
53546=>X"00",
53547=>X"00",
53548=>X"00",
53549=>X"00",
53550=>X"00",
53551=>X"00",
53552=>X"00",
53553=>X"00",
53554=>X"00",
53555=>X"00",
53556=>X"00",
53557=>X"00",
53558=>X"00",
53559=>X"00",
53560=>X"00",
53561=>X"00",
53562=>X"00",
53563=>X"00",
53564=>X"00",
53565=>X"00",
53566=>X"00",
53567=>X"00",
53568=>X"00",
53569=>X"00",
53570=>X"00",
53571=>X"00",
53572=>X"00",
53573=>X"00",
53574=>X"00",
53575=>X"00",
53576=>X"00",
53577=>X"00",
53578=>X"00",
53579=>X"00",
53580=>X"00",
53581=>X"00",
53582=>X"00",
53583=>X"00",
53584=>X"00",
53585=>X"00",
53586=>X"00",
53587=>X"00",
53588=>X"00",
53589=>X"00",
53590=>X"00",
53591=>X"00",
53592=>X"00",
53593=>X"00",
53594=>X"00",
53595=>X"00",
53596=>X"00",
53597=>X"00",
53598=>X"00",
53599=>X"00",
53600=>X"00",
53601=>X"00",
53602=>X"00",
53603=>X"00",
53604=>X"00",
53605=>X"00",
53606=>X"00",
53607=>X"00",
53608=>X"00",
53609=>X"00",
53610=>X"00",
53611=>X"00",
53612=>X"00",
53613=>X"00",
53614=>X"00",
53615=>X"00",
53616=>X"00",
53617=>X"00",
53618=>X"00",
53619=>X"00",
53620=>X"00",
53621=>X"00",
53622=>X"00",
53623=>X"00",
53624=>X"00",
53625=>X"00",
53626=>X"00",
53627=>X"00",
53628=>X"00",
53629=>X"00",
53630=>X"00",
53631=>X"00",
53632=>X"00",
53633=>X"00",
53634=>X"00",
53635=>X"00",
53636=>X"00",
53637=>X"00",
53638=>X"00",
53639=>X"00",
53640=>X"00",
53641=>X"00",
53642=>X"00",
53643=>X"00",
53644=>X"00",
53645=>X"00",
53646=>X"00",
53647=>X"00",
53648=>X"00",
53649=>X"00",
53650=>X"00",
53651=>X"00",
53652=>X"00",
53653=>X"00",
53654=>X"00",
53655=>X"00",
53656=>X"00",
53657=>X"00",
53658=>X"00",
53659=>X"00",
53660=>X"00",
53661=>X"00",
53662=>X"00",
53663=>X"00",
53664=>X"00",
53665=>X"00",
53666=>X"00",
53667=>X"00",
53668=>X"00",
53669=>X"00",
53670=>X"00",
53671=>X"00",
53672=>X"00",
53673=>X"00",
53674=>X"00",
53675=>X"00",
53676=>X"00",
53677=>X"00",
53678=>X"00",
53679=>X"00",
53680=>X"00",
53681=>X"00",
53682=>X"00",
53683=>X"00",
53684=>X"00",
53685=>X"00",
53686=>X"00",
53687=>X"00",
53688=>X"00",
53689=>X"00",
53690=>X"00",
53691=>X"00",
53692=>X"00",
53693=>X"00",
53694=>X"00",
53695=>X"00",
53696=>X"00",
53697=>X"00",
53698=>X"00",
53699=>X"00",
53700=>X"00",
53701=>X"00",
53702=>X"00",
53703=>X"00",
53704=>X"00",
53705=>X"00",
53706=>X"00",
53707=>X"00",
53708=>X"00",
53709=>X"00",
53710=>X"00",
53711=>X"00",
53712=>X"00",
53713=>X"00",
53714=>X"00",
53715=>X"00",
53716=>X"00",
53717=>X"00",
53718=>X"00",
53719=>X"00",
53720=>X"00",
53721=>X"00",
53722=>X"00",
53723=>X"00",
53724=>X"00",
53725=>X"00",
53726=>X"00",
53727=>X"00",
53728=>X"00",
53729=>X"00",
53730=>X"00",
53731=>X"00",
53732=>X"00",
53733=>X"00",
53734=>X"00",
53735=>X"00",
53736=>X"00",
53737=>X"00",
53738=>X"00",
53739=>X"00",
53740=>X"00",
53741=>X"00",
53742=>X"00",
53743=>X"00",
53744=>X"00",
53745=>X"00",
53746=>X"00",
53747=>X"00",
53748=>X"00",
53749=>X"00",
53750=>X"00",
53751=>X"00",
53752=>X"00",
53753=>X"00",
53754=>X"00",
53755=>X"00",
53756=>X"00",
53757=>X"00",
53758=>X"00",
53759=>X"00",
53760=>X"00",
53761=>X"00",
53762=>X"00",
53763=>X"00",
53764=>X"00",
53765=>X"00",
53766=>X"00",
53767=>X"00",
53768=>X"00",
53769=>X"00",
53770=>X"00",
53771=>X"00",
53772=>X"00",
53773=>X"00",
53774=>X"00",
53775=>X"00",
53776=>X"00",
53777=>X"00",
53778=>X"00",
53779=>X"00",
53780=>X"00",
53781=>X"00",
53782=>X"00",
53783=>X"00",
53784=>X"00",
53785=>X"00",
53786=>X"00",
53787=>X"00",
53788=>X"00",
53789=>X"00",
53790=>X"00",
53791=>X"00",
53792=>X"00",
53793=>X"00",
53794=>X"00",
53795=>X"00",
53796=>X"00",
53797=>X"00",
53798=>X"00",
53799=>X"00",
53800=>X"00",
53801=>X"00",
53802=>X"00",
53803=>X"00",
53804=>X"00",
53805=>X"00",
53806=>X"00",
53807=>X"00",
53808=>X"00",
53809=>X"00",
53810=>X"00",
53811=>X"00",
53812=>X"00",
53813=>X"00",
53814=>X"00",
53815=>X"00",
53816=>X"00",
53817=>X"00",
53818=>X"00",
53819=>X"00",
53820=>X"00",
53821=>X"00",
53822=>X"00",
53823=>X"00",
53824=>X"00",
53825=>X"00",
53826=>X"00",
53827=>X"00",
53828=>X"00",
53829=>X"00",
53830=>X"00",
53831=>X"00",
53832=>X"00",
53833=>X"00",
53834=>X"00",
53835=>X"00",
53836=>X"00",
53837=>X"00",
53838=>X"00",
53839=>X"00",
53840=>X"00",
53841=>X"00",
53842=>X"00",
53843=>X"00",
53844=>X"00",
53845=>X"00",
53846=>X"00",
53847=>X"00",
53848=>X"00",
53849=>X"00",
53850=>X"00",
53851=>X"00",
53852=>X"00",
53853=>X"00",
53854=>X"00",
53855=>X"00",
53856=>X"00",
53857=>X"00",
53858=>X"00",
53859=>X"00",
53860=>X"00",
53861=>X"00",
53862=>X"00",
53863=>X"00",
53864=>X"00",
53865=>X"00",
53866=>X"00",
53867=>X"00",
53868=>X"00",
53869=>X"00",
53870=>X"00",
53871=>X"00",
53872=>X"00",
53873=>X"00",
53874=>X"00",
53875=>X"00",
53876=>X"00",
53877=>X"00",
53878=>X"00",
53879=>X"00",
53880=>X"00",
53881=>X"00",
53882=>X"00",
53883=>X"00",
53884=>X"00",
53885=>X"00",
53886=>X"00",
53887=>X"00",
53888=>X"00",
53889=>X"00",
53890=>X"00",
53891=>X"00",
53892=>X"00",
53893=>X"00",
53894=>X"00",
53895=>X"00",
53896=>X"00",
53897=>X"00",
53898=>X"00",
53899=>X"00",
53900=>X"00",
53901=>X"00",
53902=>X"00",
53903=>X"00",
53904=>X"00",
53905=>X"00",
53906=>X"00",
53907=>X"00",
53908=>X"00",
53909=>X"00",
53910=>X"00",
53911=>X"00",
53912=>X"00",
53913=>X"00",
53914=>X"00",
53915=>X"00",
53916=>X"00",
53917=>X"00",
53918=>X"00",
53919=>X"00",
53920=>X"00",
53921=>X"00",
53922=>X"00",
53923=>X"00",
53924=>X"00",
53925=>X"00",
53926=>X"00",
53927=>X"00",
53928=>X"00",
53929=>X"00",
53930=>X"00",
53931=>X"00",
53932=>X"00",
53933=>X"00",
53934=>X"00",
53935=>X"00",
53936=>X"00",
53937=>X"00",
53938=>X"00",
53939=>X"00",
53940=>X"00",
53941=>X"00",
53942=>X"00",
53943=>X"00",
53944=>X"00",
53945=>X"00",
53946=>X"00",
53947=>X"00",
53948=>X"00",
53949=>X"00",
53950=>X"00",
53951=>X"00",
53952=>X"00",
53953=>X"00",
53954=>X"00",
53955=>X"00",
53956=>X"00",
53957=>X"00",
53958=>X"00",
53959=>X"00",
53960=>X"00",
53961=>X"00",
53962=>X"00",
53963=>X"00",
53964=>X"00",
53965=>X"00",
53966=>X"00",
53967=>X"00",
53968=>X"00",
53969=>X"00",
53970=>X"00",
53971=>X"00",
53972=>X"00",
53973=>X"00",
53974=>X"00",
53975=>X"00",
53976=>X"00",
53977=>X"00",
53978=>X"00",
53979=>X"00",
53980=>X"00",
53981=>X"00",
53982=>X"00",
53983=>X"00",
53984=>X"00",
53985=>X"00",
53986=>X"00",
53987=>X"00",
53988=>X"00",
53989=>X"00",
53990=>X"00",
53991=>X"00",
53992=>X"00",
53993=>X"00",
53994=>X"00",
53995=>X"00",
53996=>X"00",
53997=>X"00",
53998=>X"00",
53999=>X"00",
54000=>X"00",
54001=>X"00",
54002=>X"00",
54003=>X"00",
54004=>X"00",
54005=>X"00",
54006=>X"00",
54007=>X"00",
54008=>X"00",
54009=>X"00",
54010=>X"00",
54011=>X"00",
54012=>X"00",
54013=>X"00",
54014=>X"00",
54015=>X"00",
54016=>X"00",
54017=>X"00",
54018=>X"00",
54019=>X"00",
54020=>X"00",
54021=>X"00",
54022=>X"00",
54023=>X"00",
54024=>X"00",
54025=>X"00",
54026=>X"00",
54027=>X"00",
54028=>X"00",
54029=>X"00",
54030=>X"00",
54031=>X"00",
54032=>X"00",
54033=>X"00",
54034=>X"00",
54035=>X"00",
54036=>X"00",
54037=>X"00",
54038=>X"00",
54039=>X"00",
54040=>X"00",
54041=>X"00",
54042=>X"00",
54043=>X"00",
54044=>X"00",
54045=>X"00",
54046=>X"00",
54047=>X"00",
54048=>X"00",
54049=>X"00",
54050=>X"00",
54051=>X"00",
54052=>X"00",
54053=>X"00",
54054=>X"00",
54055=>X"00",
54056=>X"00",
54057=>X"00",
54058=>X"00",
54059=>X"00",
54060=>X"00",
54061=>X"00",
54062=>X"00",
54063=>X"00",
54064=>X"00",
54065=>X"00",
54066=>X"00",
54067=>X"00",
54068=>X"00",
54069=>X"00",
54070=>X"00",
54071=>X"00",
54072=>X"00",
54073=>X"00",
54074=>X"00",
54075=>X"00",
54076=>X"00",
54077=>X"00",
54078=>X"00",
54079=>X"00",
54080=>X"00",
54081=>X"00",
54082=>X"00",
54083=>X"00",
54084=>X"00",
54085=>X"00",
54086=>X"00",
54087=>X"00",
54088=>X"00",
54089=>X"00",
54090=>X"00",
54091=>X"00",
54092=>X"00",
54093=>X"00",
54094=>X"00",
54095=>X"00",
54096=>X"00",
54097=>X"00",
54098=>X"00",
54099=>X"00",
54100=>X"00",
54101=>X"00",
54102=>X"00",
54103=>X"00",
54104=>X"00",
54105=>X"00",
54106=>X"00",
54107=>X"00",
54108=>X"00",
54109=>X"00",
54110=>X"00",
54111=>X"00",
54112=>X"00",
54113=>X"00",
54114=>X"00",
54115=>X"00",
54116=>X"00",
54117=>X"00",
54118=>X"00",
54119=>X"00",
54120=>X"00",
54121=>X"00",
54122=>X"00",
54123=>X"00",
54124=>X"00",
54125=>X"00",
54126=>X"00",
54127=>X"00",
54128=>X"00",
54129=>X"00",
54130=>X"00",
54131=>X"00",
54132=>X"00",
54133=>X"00",
54134=>X"00",
54135=>X"00",
54136=>X"00",
54137=>X"00",
54138=>X"00",
54139=>X"00",
54140=>X"00",
54141=>X"00",
54142=>X"00",
54143=>X"00",
54144=>X"00",
54145=>X"00",
54146=>X"00",
54147=>X"00",
54148=>X"00",
54149=>X"00",
54150=>X"00",
54151=>X"00",
54152=>X"00",
54153=>X"00",
54154=>X"00",
54155=>X"00",
54156=>X"00",
54157=>X"00",
54158=>X"00",
54159=>X"00",
54160=>X"00",
54161=>X"00",
54162=>X"00",
54163=>X"00",
54164=>X"00",
54165=>X"00",
54166=>X"00",
54167=>X"00",
54168=>X"00",
54169=>X"00",
54170=>X"00",
54171=>X"00",
54172=>X"00",
54173=>X"00",
54174=>X"00",
54175=>X"00",
54176=>X"00",
54177=>X"00",
54178=>X"00",
54179=>X"00",
54180=>X"00",
54181=>X"00",
54182=>X"00",
54183=>X"00",
54184=>X"00",
54185=>X"00",
54186=>X"00",
54187=>X"00",
54188=>X"00",
54189=>X"00",
54190=>X"00",
54191=>X"00",
54192=>X"00",
54193=>X"00",
54194=>X"00",
54195=>X"00",
54196=>X"00",
54197=>X"00",
54198=>X"00",
54199=>X"00",
54200=>X"00",
54201=>X"00",
54202=>X"00",
54203=>X"00",
54204=>X"00",
54205=>X"00",
54206=>X"00",
54207=>X"00",
54208=>X"00",
54209=>X"00",
54210=>X"00",
54211=>X"00",
54212=>X"00",
54213=>X"00",
54214=>X"00",
54215=>X"00",
54216=>X"00",
54217=>X"00",
54218=>X"00",
54219=>X"00",
54220=>X"00",
54221=>X"00",
54222=>X"00",
54223=>X"00",
54224=>X"00",
54225=>X"00",
54226=>X"00",
54227=>X"00",
54228=>X"00",
54229=>X"00",
54230=>X"00",
54231=>X"00",
54232=>X"00",
54233=>X"00",
54234=>X"00",
54235=>X"00",
54236=>X"00",
54237=>X"00",
54238=>X"00",
54239=>X"00",
54240=>X"00",
54241=>X"00",
54242=>X"00",
54243=>X"00",
54244=>X"00",
54245=>X"00",
54246=>X"00",
54247=>X"00",
54248=>X"00",
54249=>X"00",
54250=>X"00",
54251=>X"00",
54252=>X"00",
54253=>X"00",
54254=>X"00",
54255=>X"00",
54256=>X"00",
54257=>X"00",
54258=>X"00",
54259=>X"00",
54260=>X"00",
54261=>X"00",
54262=>X"00",
54263=>X"00",
54264=>X"00",
54265=>X"00",
54266=>X"00",
54267=>X"00",
54268=>X"00",
54269=>X"00",
54270=>X"00",
54271=>X"00",
54272=>X"00",
54273=>X"00",
54274=>X"00",
54275=>X"00",
54276=>X"00",
54277=>X"00",
54278=>X"00",
54279=>X"00",
54280=>X"00",
54281=>X"00",
54282=>X"00",
54283=>X"00",
54284=>X"00",
54285=>X"00",
54286=>X"00",
54287=>X"00",
54288=>X"00",
54289=>X"00",
54290=>X"00",
54291=>X"00",
54292=>X"00",
54293=>X"00",
54294=>X"00",
54295=>X"00",
54296=>X"00",
54297=>X"00",
54298=>X"00",
54299=>X"00",
54300=>X"00",
54301=>X"00",
54302=>X"00",
54303=>X"00",
54304=>X"00",
54305=>X"00",
54306=>X"00",
54307=>X"00",
54308=>X"00",
54309=>X"00",
54310=>X"00",
54311=>X"00",
54312=>X"00",
54313=>X"00",
54314=>X"00",
54315=>X"00",
54316=>X"00",
54317=>X"00",
54318=>X"00",
54319=>X"00",
54320=>X"00",
54321=>X"00",
54322=>X"00",
54323=>X"00",
54324=>X"00",
54325=>X"00",
54326=>X"00",
54327=>X"00",
54328=>X"00",
54329=>X"00",
54330=>X"00",
54331=>X"00",
54332=>X"00",
54333=>X"00",
54334=>X"00",
54335=>X"00",
54336=>X"00",
54337=>X"00",
54338=>X"00",
54339=>X"00",
54340=>X"00",
54341=>X"00",
54342=>X"00",
54343=>X"00",
54344=>X"00",
54345=>X"00",
54346=>X"00",
54347=>X"00",
54348=>X"00",
54349=>X"00",
54350=>X"00",
54351=>X"00",
54352=>X"00",
54353=>X"00",
54354=>X"00",
54355=>X"00",
54356=>X"00",
54357=>X"00",
54358=>X"00",
54359=>X"00",
54360=>X"00",
54361=>X"00",
54362=>X"00",
54363=>X"00",
54364=>X"00",
54365=>X"00",
54366=>X"00",
54367=>X"00",
54368=>X"00",
54369=>X"00",
54370=>X"00",
54371=>X"00",
54372=>X"00",
54373=>X"00",
54374=>X"00",
54375=>X"00",
54376=>X"00",
54377=>X"00",
54378=>X"00",
54379=>X"00",
54380=>X"00",
54381=>X"00",
54382=>X"00",
54383=>X"00",
54384=>X"00",
54385=>X"00",
54386=>X"00",
54387=>X"00",
54388=>X"00",
54389=>X"00",
54390=>X"00",
54391=>X"00",
54392=>X"00",
54393=>X"00",
54394=>X"00",
54395=>X"00",
54396=>X"00",
54397=>X"00",
54398=>X"00",
54399=>X"00",
54400=>X"00",
54401=>X"00",
54402=>X"00",
54403=>X"00",
54404=>X"00",
54405=>X"00",
54406=>X"00",
54407=>X"00",
54408=>X"00",
54409=>X"00",
54410=>X"00",
54411=>X"00",
54412=>X"00",
54413=>X"00",
54414=>X"00",
54415=>X"00",
54416=>X"00",
54417=>X"00",
54418=>X"00",
54419=>X"00",
54420=>X"00",
54421=>X"00",
54422=>X"00",
54423=>X"00",
54424=>X"00",
54425=>X"00",
54426=>X"00",
54427=>X"00",
54428=>X"00",
54429=>X"00",
54430=>X"00",
54431=>X"00",
54432=>X"00",
54433=>X"00",
54434=>X"00",
54435=>X"00",
54436=>X"00",
54437=>X"00",
54438=>X"00",
54439=>X"00",
54440=>X"00",
54441=>X"00",
54442=>X"00",
54443=>X"00",
54444=>X"00",
54445=>X"00",
54446=>X"00",
54447=>X"00",
54448=>X"00",
54449=>X"00",
54450=>X"00",
54451=>X"00",
54452=>X"00",
54453=>X"00",
54454=>X"00",
54455=>X"00",
54456=>X"00",
54457=>X"00",
54458=>X"00",
54459=>X"00",
54460=>X"00",
54461=>X"00",
54462=>X"00",
54463=>X"00",
54464=>X"00",
54465=>X"00",
54466=>X"00",
54467=>X"00",
54468=>X"00",
54469=>X"00",
54470=>X"00",
54471=>X"00",
54472=>X"00",
54473=>X"00",
54474=>X"00",
54475=>X"00",
54476=>X"00",
54477=>X"00",
54478=>X"00",
54479=>X"00",
54480=>X"00",
54481=>X"00",
54482=>X"00",
54483=>X"00",
54484=>X"00",
54485=>X"00",
54486=>X"00",
54487=>X"00",
54488=>X"00",
54489=>X"00",
54490=>X"00",
54491=>X"00",
54492=>X"00",
54493=>X"00",
54494=>X"00",
54495=>X"00",
54496=>X"00",
54497=>X"00",
54498=>X"00",
54499=>X"00",
54500=>X"00",
54501=>X"00",
54502=>X"00",
54503=>X"00",
54504=>X"00",
54505=>X"00",
54506=>X"00",
54507=>X"00",
54508=>X"00",
54509=>X"00",
54510=>X"00",
54511=>X"00",
54512=>X"00",
54513=>X"00",
54514=>X"00",
54515=>X"00",
54516=>X"00",
54517=>X"00",
54518=>X"00",
54519=>X"00",
54520=>X"00",
54521=>X"00",
54522=>X"00",
54523=>X"00",
54524=>X"00",
54525=>X"00",
54526=>X"00",
54527=>X"00",
54528=>X"00",
54529=>X"00",
54530=>X"00",
54531=>X"00",
54532=>X"00",
54533=>X"00",
54534=>X"00",
54535=>X"00",
54536=>X"00",
54537=>X"00",
54538=>X"00",
54539=>X"00",
54540=>X"00",
54541=>X"00",
54542=>X"00",
54543=>X"00",
54544=>X"00",
54545=>X"00",
54546=>X"00",
54547=>X"00",
54548=>X"00",
54549=>X"00",
54550=>X"00",
54551=>X"00",
54552=>X"00",
54553=>X"00",
54554=>X"00",
54555=>X"00",
54556=>X"00",
54557=>X"00",
54558=>X"00",
54559=>X"00",
54560=>X"00",
54561=>X"00",
54562=>X"00",
54563=>X"00",
54564=>X"00",
54565=>X"00",
54566=>X"00",
54567=>X"00",
54568=>X"00",
54569=>X"00",
54570=>X"00",
54571=>X"00",
54572=>X"00",
54573=>X"00",
54574=>X"00",
54575=>X"00",
54576=>X"00",
54577=>X"00",
54578=>X"00",
54579=>X"00",
54580=>X"00",
54581=>X"00",
54582=>X"00",
54583=>X"00",
54584=>X"00",
54585=>X"00",
54586=>X"00",
54587=>X"00",
54588=>X"00",
54589=>X"00",
54590=>X"00",
54591=>X"00",
54592=>X"00",
54593=>X"00",
54594=>X"00",
54595=>X"00",
54596=>X"00",
54597=>X"00",
54598=>X"00",
54599=>X"00",
54600=>X"00",
54601=>X"00",
54602=>X"00",
54603=>X"00",
54604=>X"00",
54605=>X"00",
54606=>X"00",
54607=>X"00",
54608=>X"00",
54609=>X"00",
54610=>X"00",
54611=>X"00",
54612=>X"00",
54613=>X"00",
54614=>X"00",
54615=>X"00",
54616=>X"00",
54617=>X"00",
54618=>X"00",
54619=>X"00",
54620=>X"00",
54621=>X"00",
54622=>X"00",
54623=>X"00",
54624=>X"00",
54625=>X"00",
54626=>X"00",
54627=>X"00",
54628=>X"00",
54629=>X"00",
54630=>X"00",
54631=>X"00",
54632=>X"00",
54633=>X"00",
54634=>X"00",
54635=>X"00",
54636=>X"00",
54637=>X"00",
54638=>X"00",
54639=>X"00",
54640=>X"00",
54641=>X"00",
54642=>X"00",
54643=>X"00",
54644=>X"00",
54645=>X"00",
54646=>X"00",
54647=>X"00",
54648=>X"00",
54649=>X"00",
54650=>X"00",
54651=>X"00",
54652=>X"00",
54653=>X"00",
54654=>X"00",
54655=>X"00",
54656=>X"00",
54657=>X"00",
54658=>X"00",
54659=>X"00",
54660=>X"00",
54661=>X"00",
54662=>X"00",
54663=>X"00",
54664=>X"00",
54665=>X"00",
54666=>X"00",
54667=>X"00",
54668=>X"00",
54669=>X"00",
54670=>X"00",
54671=>X"00",
54672=>X"00",
54673=>X"00",
54674=>X"00",
54675=>X"00",
54676=>X"00",
54677=>X"00",
54678=>X"00",
54679=>X"00",
54680=>X"00",
54681=>X"00",
54682=>X"00",
54683=>X"00",
54684=>X"00",
54685=>X"00",
54686=>X"00",
54687=>X"00",
54688=>X"00",
54689=>X"00",
54690=>X"00",
54691=>X"00",
54692=>X"00",
54693=>X"00",
54694=>X"00",
54695=>X"00",
54696=>X"00",
54697=>X"00",
54698=>X"00",
54699=>X"00",
54700=>X"00",
54701=>X"00",
54702=>X"00",
54703=>X"00",
54704=>X"00",
54705=>X"00",
54706=>X"00",
54707=>X"00",
54708=>X"00",
54709=>X"00",
54710=>X"00",
54711=>X"00",
54712=>X"00",
54713=>X"00",
54714=>X"00",
54715=>X"00",
54716=>X"00",
54717=>X"00",
54718=>X"00",
54719=>X"00",
54720=>X"00",
54721=>X"00",
54722=>X"00",
54723=>X"00",
54724=>X"00",
54725=>X"00",
54726=>X"00",
54727=>X"00",
54728=>X"00",
54729=>X"00",
54730=>X"00",
54731=>X"00",
54732=>X"00",
54733=>X"00",
54734=>X"00",
54735=>X"00",
54736=>X"00",
54737=>X"00",
54738=>X"00",
54739=>X"00",
54740=>X"00",
54741=>X"00",
54742=>X"00",
54743=>X"00",
54744=>X"00",
54745=>X"00",
54746=>X"00",
54747=>X"00",
54748=>X"00",
54749=>X"00",
54750=>X"00",
54751=>X"00",
54752=>X"00",
54753=>X"00",
54754=>X"00",
54755=>X"00",
54756=>X"00",
54757=>X"00",
54758=>X"00",
54759=>X"00",
54760=>X"00",
54761=>X"00",
54762=>X"00",
54763=>X"00",
54764=>X"00",
54765=>X"00",
54766=>X"00",
54767=>X"00",
54768=>X"00",
54769=>X"00",
54770=>X"00",
54771=>X"00",
54772=>X"00",
54773=>X"00",
54774=>X"00",
54775=>X"00",
54776=>X"00",
54777=>X"00",
54778=>X"00",
54779=>X"00",
54780=>X"00",
54781=>X"00",
54782=>X"00",
54783=>X"00",
54784=>X"00",
54785=>X"00",
54786=>X"00",
54787=>X"00",
54788=>X"00",
54789=>X"00",
54790=>X"00",
54791=>X"00",
54792=>X"00",
54793=>X"00",
54794=>X"00",
54795=>X"00",
54796=>X"00",
54797=>X"00",
54798=>X"00",
54799=>X"00",
54800=>X"00",
54801=>X"00",
54802=>X"00",
54803=>X"00",
54804=>X"00",
54805=>X"00",
54806=>X"00",
54807=>X"00",
54808=>X"00",
54809=>X"00",
54810=>X"00",
54811=>X"00",
54812=>X"00",
54813=>X"00",
54814=>X"00",
54815=>X"00",
54816=>X"00",
54817=>X"00",
54818=>X"00",
54819=>X"00",
54820=>X"00",
54821=>X"00",
54822=>X"00",
54823=>X"00",
54824=>X"00",
54825=>X"00",
54826=>X"00",
54827=>X"00",
54828=>X"00",
54829=>X"00",
54830=>X"00",
54831=>X"00",
54832=>X"00",
54833=>X"00",
54834=>X"00",
54835=>X"00",
54836=>X"00",
54837=>X"00",
54838=>X"00",
54839=>X"00",
54840=>X"00",
54841=>X"00",
54842=>X"00",
54843=>X"00",
54844=>X"00",
54845=>X"00",
54846=>X"00",
54847=>X"00",
54848=>X"00",
54849=>X"00",
54850=>X"00",
54851=>X"00",
54852=>X"00",
54853=>X"00",
54854=>X"00",
54855=>X"00",
54856=>X"00",
54857=>X"00",
54858=>X"00",
54859=>X"00",
54860=>X"00",
54861=>X"00",
54862=>X"00",
54863=>X"00",
54864=>X"00",
54865=>X"00",
54866=>X"00",
54867=>X"00",
54868=>X"00",
54869=>X"00",
54870=>X"00",
54871=>X"00",
54872=>X"00",
54873=>X"00",
54874=>X"00",
54875=>X"00",
54876=>X"00",
54877=>X"00",
54878=>X"00",
54879=>X"00",
54880=>X"00",
54881=>X"00",
54882=>X"00",
54883=>X"00",
54884=>X"00",
54885=>X"00",
54886=>X"00",
54887=>X"00",
54888=>X"00",
54889=>X"00",
54890=>X"00",
54891=>X"00",
54892=>X"00",
54893=>X"00",
54894=>X"00",
54895=>X"00",
54896=>X"00",
54897=>X"00",
54898=>X"00",
54899=>X"00",
54900=>X"00",
54901=>X"00",
54902=>X"00",
54903=>X"00",
54904=>X"00",
54905=>X"00",
54906=>X"00",
54907=>X"00",
54908=>X"00",
54909=>X"00",
54910=>X"00",
54911=>X"00",
54912=>X"00",
54913=>X"00",
54914=>X"00",
54915=>X"00",
54916=>X"00",
54917=>X"00",
54918=>X"00",
54919=>X"00",
54920=>X"00",
54921=>X"00",
54922=>X"00",
54923=>X"00",
54924=>X"00",
54925=>X"00",
54926=>X"00",
54927=>X"00",
54928=>X"00",
54929=>X"00",
54930=>X"00",
54931=>X"00",
54932=>X"00",
54933=>X"00",
54934=>X"00",
54935=>X"00",
54936=>X"00",
54937=>X"00",
54938=>X"00",
54939=>X"00",
54940=>X"00",
54941=>X"00",
54942=>X"00",
54943=>X"00",
54944=>X"00",
54945=>X"00",
54946=>X"00",
54947=>X"00",
54948=>X"00",
54949=>X"00",
54950=>X"00",
54951=>X"00",
54952=>X"00",
54953=>X"00",
54954=>X"00",
54955=>X"00",
54956=>X"00",
54957=>X"00",
54958=>X"00",
54959=>X"00",
54960=>X"00",
54961=>X"00",
54962=>X"00",
54963=>X"00",
54964=>X"00",
54965=>X"00",
54966=>X"00",
54967=>X"00",
54968=>X"00",
54969=>X"00",
54970=>X"00",
54971=>X"00",
54972=>X"00",
54973=>X"00",
54974=>X"00",
54975=>X"00",
54976=>X"00",
54977=>X"00",
54978=>X"00",
54979=>X"00",
54980=>X"00",
54981=>X"00",
54982=>X"00",
54983=>X"00",
54984=>X"00",
54985=>X"00",
54986=>X"00",
54987=>X"00",
54988=>X"00",
54989=>X"00",
54990=>X"00",
54991=>X"00",
54992=>X"00",
54993=>X"00",
54994=>X"00",
54995=>X"00",
54996=>X"00",
54997=>X"00",
54998=>X"00",
54999=>X"00",
55000=>X"00",
55001=>X"00",
55002=>X"00",
55003=>X"00",
55004=>X"00",
55005=>X"00",
55006=>X"00",
55007=>X"00",
55008=>X"00",
55009=>X"00",
55010=>X"00",
55011=>X"00",
55012=>X"00",
55013=>X"00",
55014=>X"00",
55015=>X"00",
55016=>X"00",
55017=>X"00",
55018=>X"00",
55019=>X"00",
55020=>X"00",
55021=>X"00",
55022=>X"00",
55023=>X"00",
55024=>X"00",
55025=>X"00",
55026=>X"00",
55027=>X"00",
55028=>X"00",
55029=>X"00",
55030=>X"00",
55031=>X"00",
55032=>X"00",
55033=>X"00",
55034=>X"00",
55035=>X"00",
55036=>X"00",
55037=>X"00",
55038=>X"00",
55039=>X"00",
55040=>X"00",
55041=>X"00",
55042=>X"00",
55043=>X"00",
55044=>X"00",
55045=>X"00",
55046=>X"00",
55047=>X"00",
55048=>X"00",
55049=>X"00",
55050=>X"00",
55051=>X"00",
55052=>X"00",
55053=>X"00",
55054=>X"00",
55055=>X"00",
55056=>X"00",
55057=>X"00",
55058=>X"00",
55059=>X"00",
55060=>X"00",
55061=>X"00",
55062=>X"00",
55063=>X"00",
55064=>X"00",
55065=>X"00",
55066=>X"00",
55067=>X"00",
55068=>X"00",
55069=>X"00",
55070=>X"00",
55071=>X"00",
55072=>X"00",
55073=>X"00",
55074=>X"00",
55075=>X"00",
55076=>X"00",
55077=>X"00",
55078=>X"00",
55079=>X"00",
55080=>X"00",
55081=>X"00",
55082=>X"00",
55083=>X"00",
55084=>X"00",
55085=>X"00",
55086=>X"00",
55087=>X"00",
55088=>X"00",
55089=>X"00",
55090=>X"00",
55091=>X"00",
55092=>X"00",
55093=>X"00",
55094=>X"00",
55095=>X"00",
55096=>X"00",
55097=>X"00",
55098=>X"00",
55099=>X"00",
55100=>X"00",
55101=>X"00",
55102=>X"00",
55103=>X"00",
55104=>X"00",
55105=>X"00",
55106=>X"00",
55107=>X"00",
55108=>X"00",
55109=>X"00",
55110=>X"00",
55111=>X"00",
55112=>X"00",
55113=>X"00",
55114=>X"00",
55115=>X"00",
55116=>X"00",
55117=>X"00",
55118=>X"00",
55119=>X"00",
55120=>X"00",
55121=>X"00",
55122=>X"00",
55123=>X"00",
55124=>X"00",
55125=>X"00",
55126=>X"00",
55127=>X"00",
55128=>X"00",
55129=>X"00",
55130=>X"00",
55131=>X"00",
55132=>X"00",
55133=>X"00",
55134=>X"00",
55135=>X"00",
55136=>X"00",
55137=>X"00",
55138=>X"00",
55139=>X"00",
55140=>X"00",
55141=>X"00",
55142=>X"00",
55143=>X"00",
55144=>X"00",
55145=>X"00",
55146=>X"00",
55147=>X"00",
55148=>X"00",
55149=>X"00",
55150=>X"00",
55151=>X"00",
55152=>X"00",
55153=>X"00",
55154=>X"00",
55155=>X"00",
55156=>X"00",
55157=>X"00",
55158=>X"00",
55159=>X"00",
55160=>X"00",
55161=>X"00",
55162=>X"00",
55163=>X"00",
55164=>X"00",
55165=>X"00",
55166=>X"00",
55167=>X"00",
55168=>X"00",
55169=>X"00",
55170=>X"00",
55171=>X"00",
55172=>X"00",
55173=>X"00",
55174=>X"00",
55175=>X"00",
55176=>X"00",
55177=>X"00",
55178=>X"00",
55179=>X"00",
55180=>X"00",
55181=>X"00",
55182=>X"00",
55183=>X"00",
55184=>X"00",
55185=>X"00",
55186=>X"00",
55187=>X"00",
55188=>X"00",
55189=>X"00",
55190=>X"00",
55191=>X"00",
55192=>X"00",
55193=>X"00",
55194=>X"00",
55195=>X"00",
55196=>X"00",
55197=>X"00",
55198=>X"00",
55199=>X"00",
55200=>X"00",
55201=>X"00",
55202=>X"00",
55203=>X"00",
55204=>X"00",
55205=>X"00",
55206=>X"00",
55207=>X"00",
55208=>X"00",
55209=>X"00",
55210=>X"00",
55211=>X"00",
55212=>X"00",
55213=>X"00",
55214=>X"00",
55215=>X"00",
55216=>X"00",
55217=>X"00",
55218=>X"00",
55219=>X"00",
55220=>X"00",
55221=>X"00",
55222=>X"00",
55223=>X"00",
55224=>X"00",
55225=>X"00",
55226=>X"00",
55227=>X"00",
55228=>X"00",
55229=>X"00",
55230=>X"00",
55231=>X"00",
55232=>X"00",
55233=>X"00",
55234=>X"00",
55235=>X"00",
55236=>X"00",
55237=>X"00",
55238=>X"00",
55239=>X"00",
55240=>X"00",
55241=>X"00",
55242=>X"00",
55243=>X"00",
55244=>X"00",
55245=>X"00",
55246=>X"00",
55247=>X"00",
55248=>X"00",
55249=>X"00",
55250=>X"00",
55251=>X"00",
55252=>X"00",
55253=>X"00",
55254=>X"00",
55255=>X"00",
55256=>X"00",
55257=>X"00",
55258=>X"00",
55259=>X"00",
55260=>X"00",
55261=>X"00",
55262=>X"00",
55263=>X"00",
55264=>X"00",
55265=>X"00",
55266=>X"00",
55267=>X"00",
55268=>X"00",
55269=>X"00",
55270=>X"00",
55271=>X"00",
55272=>X"00",
55273=>X"00",
55274=>X"00",
55275=>X"00",
55276=>X"00",
55277=>X"00",
55278=>X"00",
55279=>X"00",
55280=>X"00",
55281=>X"00",
55282=>X"00",
55283=>X"00",
55284=>X"00",
55285=>X"00",
55286=>X"00",
55287=>X"00",
55288=>X"00",
55289=>X"00",
55290=>X"00",
55291=>X"00",
55292=>X"00",
55293=>X"00",
55294=>X"00",
55295=>X"00",
55296=>X"00",
55297=>X"00",
55298=>X"00",
55299=>X"00",
55300=>X"00",
55301=>X"00",
55302=>X"00",
55303=>X"00",
55304=>X"00",
55305=>X"00",
55306=>X"00",
55307=>X"00",
55308=>X"00",
55309=>X"00",
55310=>X"00",
55311=>X"00",
55312=>X"00",
55313=>X"00",
55314=>X"00",
55315=>X"00",
55316=>X"00",
55317=>X"00",
55318=>X"00",
55319=>X"00",
55320=>X"00",
55321=>X"00",
55322=>X"00",
55323=>X"00",
55324=>X"00",
55325=>X"00",
55326=>X"00",
55327=>X"00",
55328=>X"00",
55329=>X"00",
55330=>X"00",
55331=>X"00",
55332=>X"00",
55333=>X"00",
55334=>X"00",
55335=>X"00",
55336=>X"00",
55337=>X"00",
55338=>X"00",
55339=>X"00",
55340=>X"00",
55341=>X"00",
55342=>X"00",
55343=>X"00",
55344=>X"00",
55345=>X"00",
55346=>X"00",
55347=>X"00",
55348=>X"00",
55349=>X"00",
55350=>X"00",
55351=>X"00",
55352=>X"00",
55353=>X"00",
55354=>X"00",
55355=>X"00",
55356=>X"00",
55357=>X"00",
55358=>X"00",
55359=>X"00",
55360=>X"00",
55361=>X"00",
55362=>X"00",
55363=>X"00",
55364=>X"00",
55365=>X"00",
55366=>X"00",
55367=>X"00",
55368=>X"00",
55369=>X"00",
55370=>X"00",
55371=>X"00",
55372=>X"00",
55373=>X"00",
55374=>X"00",
55375=>X"00",
55376=>X"00",
55377=>X"00",
55378=>X"00",
55379=>X"00",
55380=>X"00",
55381=>X"00",
55382=>X"00",
55383=>X"00",
55384=>X"00",
55385=>X"00",
55386=>X"00",
55387=>X"00",
55388=>X"00",
55389=>X"00",
55390=>X"00",
55391=>X"00",
55392=>X"00",
55393=>X"00",
55394=>X"00",
55395=>X"00",
55396=>X"00",
55397=>X"00",
55398=>X"00",
55399=>X"00",
55400=>X"00",
55401=>X"00",
55402=>X"00",
55403=>X"00",
55404=>X"00",
55405=>X"00",
55406=>X"00",
55407=>X"00",
55408=>X"00",
55409=>X"00",
55410=>X"00",
55411=>X"00",
55412=>X"00",
55413=>X"00",
55414=>X"00",
55415=>X"00",
55416=>X"00",
55417=>X"00",
55418=>X"00",
55419=>X"00",
55420=>X"00",
55421=>X"00",
55422=>X"00",
55423=>X"00",
55424=>X"00",
55425=>X"00",
55426=>X"00",
55427=>X"00",
55428=>X"00",
55429=>X"00",
55430=>X"00",
55431=>X"00",
55432=>X"00",
55433=>X"00",
55434=>X"00",
55435=>X"00",
55436=>X"00",
55437=>X"00",
55438=>X"00",
55439=>X"00",
55440=>X"00",
55441=>X"00",
55442=>X"00",
55443=>X"00",
55444=>X"00",
55445=>X"00",
55446=>X"00",
55447=>X"00",
55448=>X"00",
55449=>X"00",
55450=>X"00",
55451=>X"00",
55452=>X"00",
55453=>X"00",
55454=>X"00",
55455=>X"00",
55456=>X"00",
55457=>X"00",
55458=>X"00",
55459=>X"00",
55460=>X"00",
55461=>X"00",
55462=>X"00",
55463=>X"00",
55464=>X"00",
55465=>X"00",
55466=>X"00",
55467=>X"00",
55468=>X"00",
55469=>X"00",
55470=>X"00",
55471=>X"00",
55472=>X"00",
55473=>X"00",
55474=>X"00",
55475=>X"00",
55476=>X"00",
55477=>X"00",
55478=>X"00",
55479=>X"00",
55480=>X"00",
55481=>X"00",
55482=>X"00",
55483=>X"00",
55484=>X"00",
55485=>X"00",
55486=>X"00",
55487=>X"00",
55488=>X"00",
55489=>X"00",
55490=>X"00",
55491=>X"00",
55492=>X"00",
55493=>X"00",
55494=>X"00",
55495=>X"00",
55496=>X"00",
55497=>X"00",
55498=>X"00",
55499=>X"00",
55500=>X"00",
55501=>X"00",
55502=>X"00",
55503=>X"00",
55504=>X"00",
55505=>X"00",
55506=>X"00",
55507=>X"00",
55508=>X"00",
55509=>X"00",
55510=>X"00",
55511=>X"00",
55512=>X"00",
55513=>X"00",
55514=>X"00",
55515=>X"00",
55516=>X"00",
55517=>X"00",
55518=>X"00",
55519=>X"00",
55520=>X"00",
55521=>X"00",
55522=>X"00",
55523=>X"00",
55524=>X"00",
55525=>X"00",
55526=>X"00",
55527=>X"00",
55528=>X"00",
55529=>X"00",
55530=>X"00",
55531=>X"00",
55532=>X"00",
55533=>X"00",
55534=>X"00",
55535=>X"00",
55536=>X"00",
55537=>X"00",
55538=>X"00",
55539=>X"00",
55540=>X"00",
55541=>X"00",
55542=>X"00",
55543=>X"00",
55544=>X"00",
55545=>X"00",
55546=>X"00",
55547=>X"00",
55548=>X"00",
55549=>X"00",
55550=>X"00",
55551=>X"00",
55552=>X"00",
55553=>X"00",
55554=>X"00",
55555=>X"00",
55556=>X"00",
55557=>X"00",
55558=>X"00",
55559=>X"00",
55560=>X"00",
55561=>X"00",
55562=>X"00",
55563=>X"00",
55564=>X"00",
55565=>X"00",
55566=>X"00",
55567=>X"00",
55568=>X"00",
55569=>X"00",
55570=>X"00",
55571=>X"00",
55572=>X"00",
55573=>X"00",
55574=>X"00",
55575=>X"00",
55576=>X"00",
55577=>X"00",
55578=>X"00",
55579=>X"00",
55580=>X"00",
55581=>X"00",
55582=>X"00",
55583=>X"00",
55584=>X"00",
55585=>X"00",
55586=>X"00",
55587=>X"00",
55588=>X"00",
55589=>X"00",
55590=>X"00",
55591=>X"00",
55592=>X"00",
55593=>X"00",
55594=>X"00",
55595=>X"00",
55596=>X"00",
55597=>X"00",
55598=>X"00",
55599=>X"00",
55600=>X"00",
55601=>X"00",
55602=>X"00",
55603=>X"00",
55604=>X"00",
55605=>X"00",
55606=>X"00",
55607=>X"00",
55608=>X"00",
55609=>X"00",
55610=>X"00",
55611=>X"00",
55612=>X"00",
55613=>X"00",
55614=>X"00",
55615=>X"00",
55616=>X"00",
55617=>X"00",
55618=>X"00",
55619=>X"00",
55620=>X"00",
55621=>X"00",
55622=>X"00",
55623=>X"00",
55624=>X"00",
55625=>X"00",
55626=>X"00",
55627=>X"00",
55628=>X"00",
55629=>X"00",
55630=>X"00",
55631=>X"00",
55632=>X"00",
55633=>X"00",
55634=>X"00",
55635=>X"00",
55636=>X"00",
55637=>X"00",
55638=>X"00",
55639=>X"00",
55640=>X"00",
55641=>X"00",
55642=>X"00",
55643=>X"00",
55644=>X"00",
55645=>X"00",
55646=>X"00",
55647=>X"00",
55648=>X"00",
55649=>X"00",
55650=>X"00",
55651=>X"00",
55652=>X"00",
55653=>X"00",
55654=>X"00",
55655=>X"00",
55656=>X"00",
55657=>X"00",
55658=>X"00",
55659=>X"00",
55660=>X"00",
55661=>X"00",
55662=>X"00",
55663=>X"00",
55664=>X"00",
55665=>X"00",
55666=>X"00",
55667=>X"00",
55668=>X"00",
55669=>X"00",
55670=>X"00",
55671=>X"00",
55672=>X"00",
55673=>X"00",
55674=>X"00",
55675=>X"00",
55676=>X"00",
55677=>X"00",
55678=>X"00",
55679=>X"00",
55680=>X"00",
55681=>X"00",
55682=>X"00",
55683=>X"00",
55684=>X"00",
55685=>X"00",
55686=>X"00",
55687=>X"00",
55688=>X"00",
55689=>X"00",
55690=>X"00",
55691=>X"00",
55692=>X"00",
55693=>X"00",
55694=>X"00",
55695=>X"00",
55696=>X"00",
55697=>X"00",
55698=>X"00",
55699=>X"00",
55700=>X"00",
55701=>X"00",
55702=>X"00",
55703=>X"00",
55704=>X"00",
55705=>X"00",
55706=>X"00",
55707=>X"00",
55708=>X"00",
55709=>X"00",
55710=>X"00",
55711=>X"00",
55712=>X"00",
55713=>X"00",
55714=>X"00",
55715=>X"00",
55716=>X"00",
55717=>X"00",
55718=>X"00",
55719=>X"00",
55720=>X"00",
55721=>X"00",
55722=>X"00",
55723=>X"00",
55724=>X"00",
55725=>X"00",
55726=>X"00",
55727=>X"00",
55728=>X"00",
55729=>X"00",
55730=>X"00",
55731=>X"00",
55732=>X"00",
55733=>X"00",
55734=>X"00",
55735=>X"00",
55736=>X"00",
55737=>X"00",
55738=>X"00",
55739=>X"00",
55740=>X"00",
55741=>X"00",
55742=>X"00",
55743=>X"00",
55744=>X"00",
55745=>X"00",
55746=>X"00",
55747=>X"00",
55748=>X"00",
55749=>X"00",
55750=>X"00",
55751=>X"00",
55752=>X"00",
55753=>X"00",
55754=>X"00",
55755=>X"00",
55756=>X"00",
55757=>X"00",
55758=>X"00",
55759=>X"00",
55760=>X"00",
55761=>X"00",
55762=>X"00",
55763=>X"00",
55764=>X"00",
55765=>X"00",
55766=>X"00",
55767=>X"00",
55768=>X"00",
55769=>X"00",
55770=>X"00",
55771=>X"00",
55772=>X"00",
55773=>X"00",
55774=>X"00",
55775=>X"00",
55776=>X"00",
55777=>X"00",
55778=>X"00",
55779=>X"00",
55780=>X"00",
55781=>X"00",
55782=>X"00",
55783=>X"00",
55784=>X"00",
55785=>X"00",
55786=>X"00",
55787=>X"00",
55788=>X"00",
55789=>X"00",
55790=>X"00",
55791=>X"00",
55792=>X"00",
55793=>X"00",
55794=>X"00",
55795=>X"00",
55796=>X"00",
55797=>X"00",
55798=>X"00",
55799=>X"00",
55800=>X"00",
55801=>X"00",
55802=>X"00",
55803=>X"00",
55804=>X"00",
55805=>X"00",
55806=>X"00",
55807=>X"00",
55808=>X"00",
55809=>X"00",
55810=>X"00",
55811=>X"00",
55812=>X"00",
55813=>X"00",
55814=>X"00",
55815=>X"00",
55816=>X"00",
55817=>X"00",
55818=>X"00",
55819=>X"00",
55820=>X"00",
55821=>X"00",
55822=>X"00",
55823=>X"00",
55824=>X"00",
55825=>X"00",
55826=>X"00",
55827=>X"00",
55828=>X"00",
55829=>X"00",
55830=>X"00",
55831=>X"00",
55832=>X"00",
55833=>X"00",
55834=>X"00",
55835=>X"00",
55836=>X"00",
55837=>X"00",
55838=>X"00",
55839=>X"00",
55840=>X"00",
55841=>X"00",
55842=>X"00",
55843=>X"00",
55844=>X"00",
55845=>X"00",
55846=>X"00",
55847=>X"00",
55848=>X"00",
55849=>X"00",
55850=>X"00",
55851=>X"00",
55852=>X"00",
55853=>X"00",
55854=>X"00",
55855=>X"00",
55856=>X"00",
55857=>X"00",
55858=>X"00",
55859=>X"00",
55860=>X"00",
55861=>X"00",
55862=>X"00",
55863=>X"00",
55864=>X"00",
55865=>X"00",
55866=>X"00",
55867=>X"00",
55868=>X"00",
55869=>X"00",
55870=>X"00",
55871=>X"00",
55872=>X"00",
55873=>X"00",
55874=>X"00",
55875=>X"00",
55876=>X"00",
55877=>X"00",
55878=>X"00",
55879=>X"00",
55880=>X"00",
55881=>X"00",
55882=>X"00",
55883=>X"00",
55884=>X"00",
55885=>X"00",
55886=>X"00",
55887=>X"00",
55888=>X"00",
55889=>X"00",
55890=>X"00",
55891=>X"00",
55892=>X"00",
55893=>X"00",
55894=>X"00",
55895=>X"00",
55896=>X"00",
55897=>X"00",
55898=>X"00",
55899=>X"00",
55900=>X"00",
55901=>X"00",
55902=>X"00",
55903=>X"00",
55904=>X"00",
55905=>X"00",
55906=>X"00",
55907=>X"00",
55908=>X"00",
55909=>X"00",
55910=>X"00",
55911=>X"00",
55912=>X"00",
55913=>X"00",
55914=>X"00",
55915=>X"00",
55916=>X"00",
55917=>X"00",
55918=>X"00",
55919=>X"00",
55920=>X"00",
55921=>X"00",
55922=>X"00",
55923=>X"00",
55924=>X"00",
55925=>X"00",
55926=>X"00",
55927=>X"00",
55928=>X"00",
55929=>X"00",
55930=>X"00",
55931=>X"00",
55932=>X"00",
55933=>X"00",
55934=>X"00",
55935=>X"00",
55936=>X"00",
55937=>X"00",
55938=>X"00",
55939=>X"00",
55940=>X"00",
55941=>X"00",
55942=>X"00",
55943=>X"00",
55944=>X"00",
55945=>X"00",
55946=>X"00",
55947=>X"00",
55948=>X"00",
55949=>X"00",
55950=>X"00",
55951=>X"00",
55952=>X"00",
55953=>X"00",
55954=>X"00",
55955=>X"00",
55956=>X"00",
55957=>X"00",
55958=>X"00",
55959=>X"00",
55960=>X"00",
55961=>X"00",
55962=>X"00",
55963=>X"00",
55964=>X"00",
55965=>X"00",
55966=>X"00",
55967=>X"00",
55968=>X"00",
55969=>X"00",
55970=>X"00",
55971=>X"00",
55972=>X"00",
55973=>X"00",
55974=>X"00",
55975=>X"00",
55976=>X"00",
55977=>X"00",
55978=>X"00",
55979=>X"00",
55980=>X"00",
55981=>X"00",
55982=>X"00",
55983=>X"00",
55984=>X"00",
55985=>X"00",
55986=>X"00",
55987=>X"00",
55988=>X"00",
55989=>X"00",
55990=>X"00",
55991=>X"00",
55992=>X"00",
55993=>X"00",
55994=>X"00",
55995=>X"00",
55996=>X"00",
55997=>X"00",
55998=>X"00",
55999=>X"00",
56000=>X"00",
56001=>X"00",
56002=>X"00",
56003=>X"00",
56004=>X"00",
56005=>X"00",
56006=>X"00",
56007=>X"00",
56008=>X"00",
56009=>X"00",
56010=>X"00",
56011=>X"00",
56012=>X"00",
56013=>X"00",
56014=>X"00",
56015=>X"00",
56016=>X"00",
56017=>X"00",
56018=>X"00",
56019=>X"00",
56020=>X"00",
56021=>X"00",
56022=>X"00",
56023=>X"00",
56024=>X"00",
56025=>X"00",
56026=>X"00",
56027=>X"00",
56028=>X"00",
56029=>X"00",
56030=>X"00",
56031=>X"00",
56032=>X"00",
56033=>X"00",
56034=>X"00",
56035=>X"00",
56036=>X"00",
56037=>X"00",
56038=>X"00",
56039=>X"00",
56040=>X"00",
56041=>X"00",
56042=>X"00",
56043=>X"00",
56044=>X"00",
56045=>X"00",
56046=>X"00",
56047=>X"00",
56048=>X"00",
56049=>X"00",
56050=>X"00",
56051=>X"00",
56052=>X"00",
56053=>X"00",
56054=>X"00",
56055=>X"00",
56056=>X"00",
56057=>X"00",
56058=>X"00",
56059=>X"00",
56060=>X"00",
56061=>X"00",
56062=>X"00",
56063=>X"00",
56064=>X"00",
56065=>X"00",
56066=>X"00",
56067=>X"00",
56068=>X"00",
56069=>X"00",
56070=>X"00",
56071=>X"00",
56072=>X"00",
56073=>X"00",
56074=>X"00",
56075=>X"00",
56076=>X"00",
56077=>X"00",
56078=>X"00",
56079=>X"00",
56080=>X"00",
56081=>X"00",
56082=>X"00",
56083=>X"00",
56084=>X"00",
56085=>X"00",
56086=>X"00",
56087=>X"00",
56088=>X"00",
56089=>X"00",
56090=>X"00",
56091=>X"00",
56092=>X"00",
56093=>X"00",
56094=>X"00",
56095=>X"00",
56096=>X"00",
56097=>X"00",
56098=>X"00",
56099=>X"00",
56100=>X"00",
56101=>X"00",
56102=>X"00",
56103=>X"00",
56104=>X"00",
56105=>X"00",
56106=>X"00",
56107=>X"00",
56108=>X"00",
56109=>X"00",
56110=>X"00",
56111=>X"00",
56112=>X"00",
56113=>X"00",
56114=>X"00",
56115=>X"00",
56116=>X"00",
56117=>X"00",
56118=>X"00",
56119=>X"00",
56120=>X"00",
56121=>X"00",
56122=>X"00",
56123=>X"00",
56124=>X"00",
56125=>X"00",
56126=>X"00",
56127=>X"00",
56128=>X"00",
56129=>X"00",
56130=>X"00",
56131=>X"00",
56132=>X"00",
56133=>X"00",
56134=>X"00",
56135=>X"00",
56136=>X"00",
56137=>X"00",
56138=>X"00",
56139=>X"00",
56140=>X"00",
56141=>X"00",
56142=>X"00",
56143=>X"00",
56144=>X"00",
56145=>X"00",
56146=>X"00",
56147=>X"00",
56148=>X"00",
56149=>X"00",
56150=>X"00",
56151=>X"00",
56152=>X"00",
56153=>X"00",
56154=>X"00",
56155=>X"00",
56156=>X"00",
56157=>X"00",
56158=>X"00",
56159=>X"00",
56160=>X"00",
56161=>X"00",
56162=>X"00",
56163=>X"00",
56164=>X"00",
56165=>X"00",
56166=>X"00",
56167=>X"00",
56168=>X"00",
56169=>X"00",
56170=>X"00",
56171=>X"00",
56172=>X"00",
56173=>X"00",
56174=>X"00",
56175=>X"00",
56176=>X"00",
56177=>X"00",
56178=>X"00",
56179=>X"00",
56180=>X"00",
56181=>X"00",
56182=>X"00",
56183=>X"00",
56184=>X"00",
56185=>X"00",
56186=>X"00",
56187=>X"00",
56188=>X"00",
56189=>X"00",
56190=>X"00",
56191=>X"00",
56192=>X"00",
56193=>X"00",
56194=>X"00",
56195=>X"00",
56196=>X"00",
56197=>X"00",
56198=>X"00",
56199=>X"00",
56200=>X"00",
56201=>X"00",
56202=>X"00",
56203=>X"00",
56204=>X"00",
56205=>X"00",
56206=>X"00",
56207=>X"00",
56208=>X"00",
56209=>X"00",
56210=>X"00",
56211=>X"00",
56212=>X"00",
56213=>X"00",
56214=>X"00",
56215=>X"00",
56216=>X"00",
56217=>X"00",
56218=>X"00",
56219=>X"00",
56220=>X"00",
56221=>X"00",
56222=>X"00",
56223=>X"00",
56224=>X"00",
56225=>X"00",
56226=>X"00",
56227=>X"00",
56228=>X"00",
56229=>X"00",
56230=>X"00",
56231=>X"00",
56232=>X"00",
56233=>X"00",
56234=>X"00",
56235=>X"00",
56236=>X"00",
56237=>X"00",
56238=>X"00",
56239=>X"00",
56240=>X"00",
56241=>X"00",
56242=>X"00",
56243=>X"00",
56244=>X"00",
56245=>X"00",
56246=>X"00",
56247=>X"00",
56248=>X"00",
56249=>X"00",
56250=>X"00",
56251=>X"00",
56252=>X"00",
56253=>X"00",
56254=>X"00",
56255=>X"00",
56256=>X"00",
56257=>X"00",
56258=>X"00",
56259=>X"00",
56260=>X"00",
56261=>X"00",
56262=>X"00",
56263=>X"00",
56264=>X"00",
56265=>X"00",
56266=>X"00",
56267=>X"00",
56268=>X"00",
56269=>X"00",
56270=>X"00",
56271=>X"00",
56272=>X"00",
56273=>X"00",
56274=>X"00",
56275=>X"00",
56276=>X"00",
56277=>X"00",
56278=>X"00",
56279=>X"00",
56280=>X"00",
56281=>X"00",
56282=>X"00",
56283=>X"00",
56284=>X"00",
56285=>X"00",
56286=>X"00",
56287=>X"00",
56288=>X"00",
56289=>X"00",
56290=>X"00",
56291=>X"00",
56292=>X"00",
56293=>X"00",
56294=>X"00",
56295=>X"00",
56296=>X"00",
56297=>X"00",
56298=>X"00",
56299=>X"00",
56300=>X"00",
56301=>X"00",
56302=>X"00",
56303=>X"00",
56304=>X"00",
56305=>X"00",
56306=>X"00",
56307=>X"00",
56308=>X"00",
56309=>X"00",
56310=>X"00",
56311=>X"00",
56312=>X"00",
56313=>X"00",
56314=>X"00",
56315=>X"00",
56316=>X"00",
56317=>X"00",
56318=>X"00",
56319=>X"00",
56320=>X"00",
56321=>X"00",
56322=>X"00",
56323=>X"00",
56324=>X"00",
56325=>X"00",
56326=>X"00",
56327=>X"00",
56328=>X"00",
56329=>X"00",
56330=>X"00",
56331=>X"00",
56332=>X"00",
56333=>X"00",
56334=>X"00",
56335=>X"00",
56336=>X"00",
56337=>X"00",
56338=>X"00",
56339=>X"00",
56340=>X"00",
56341=>X"00",
56342=>X"00",
56343=>X"00",
56344=>X"00",
56345=>X"00",
56346=>X"00",
56347=>X"00",
56348=>X"00",
56349=>X"00",
56350=>X"00",
56351=>X"00",
56352=>X"00",
56353=>X"00",
56354=>X"00",
56355=>X"00",
56356=>X"00",
56357=>X"00",
56358=>X"00",
56359=>X"00",
56360=>X"00",
56361=>X"00",
56362=>X"00",
56363=>X"00",
56364=>X"00",
56365=>X"00",
56366=>X"00",
56367=>X"00",
56368=>X"00",
56369=>X"00",
56370=>X"00",
56371=>X"00",
56372=>X"00",
56373=>X"00",
56374=>X"00",
56375=>X"00",
56376=>X"00",
56377=>X"00",
56378=>X"00",
56379=>X"00",
56380=>X"00",
56381=>X"00",
56382=>X"00",
56383=>X"00",
56384=>X"00",
56385=>X"00",
56386=>X"00",
56387=>X"00",
56388=>X"00",
56389=>X"00",
56390=>X"00",
56391=>X"00",
56392=>X"00",
56393=>X"00",
56394=>X"00",
56395=>X"00",
56396=>X"00",
56397=>X"00",
56398=>X"00",
56399=>X"00",
56400=>X"00",
56401=>X"00",
56402=>X"00",
56403=>X"00",
56404=>X"00",
56405=>X"00",
56406=>X"00",
56407=>X"00",
56408=>X"00",
56409=>X"00",
56410=>X"00",
56411=>X"00",
56412=>X"00",
56413=>X"00",
56414=>X"00",
56415=>X"00",
56416=>X"00",
56417=>X"00",
56418=>X"00",
56419=>X"00",
56420=>X"00",
56421=>X"00",
56422=>X"00",
56423=>X"00",
56424=>X"00",
56425=>X"00",
56426=>X"00",
56427=>X"00",
56428=>X"00",
56429=>X"00",
56430=>X"00",
56431=>X"00",
56432=>X"00",
56433=>X"00",
56434=>X"00",
56435=>X"00",
56436=>X"00",
56437=>X"00",
56438=>X"00",
56439=>X"00",
56440=>X"00",
56441=>X"00",
56442=>X"00",
56443=>X"00",
56444=>X"00",
56445=>X"00",
56446=>X"00",
56447=>X"00",
56448=>X"00",
56449=>X"00",
56450=>X"00",
56451=>X"00",
56452=>X"00",
56453=>X"00",
56454=>X"00",
56455=>X"00",
56456=>X"00",
56457=>X"00",
56458=>X"00",
56459=>X"00",
56460=>X"00",
56461=>X"00",
56462=>X"00",
56463=>X"00",
56464=>X"00",
56465=>X"00",
56466=>X"00",
56467=>X"00",
56468=>X"00",
56469=>X"00",
56470=>X"00",
56471=>X"00",
56472=>X"00",
56473=>X"00",
56474=>X"00",
56475=>X"00",
56476=>X"00",
56477=>X"00",
56478=>X"00",
56479=>X"00",
56480=>X"00",
56481=>X"00",
56482=>X"00",
56483=>X"00",
56484=>X"00",
56485=>X"00",
56486=>X"00",
56487=>X"00",
56488=>X"00",
56489=>X"00",
56490=>X"00",
56491=>X"00",
56492=>X"00",
56493=>X"00",
56494=>X"00",
56495=>X"00",
56496=>X"00",
56497=>X"00",
56498=>X"00",
56499=>X"00",
56500=>X"00",
56501=>X"00",
56502=>X"00",
56503=>X"00",
56504=>X"00",
56505=>X"00",
56506=>X"00",
56507=>X"00",
56508=>X"00",
56509=>X"00",
56510=>X"00",
56511=>X"00",
56512=>X"00",
56513=>X"00",
56514=>X"00",
56515=>X"00",
56516=>X"00",
56517=>X"00",
56518=>X"00",
56519=>X"00",
56520=>X"00",
56521=>X"00",
56522=>X"00",
56523=>X"00",
56524=>X"00",
56525=>X"00",
56526=>X"00",
56527=>X"00",
56528=>X"00",
56529=>X"00",
56530=>X"00",
56531=>X"00",
56532=>X"00",
56533=>X"00",
56534=>X"00",
56535=>X"00",
56536=>X"00",
56537=>X"00",
56538=>X"00",
56539=>X"00",
56540=>X"00",
56541=>X"00",
56542=>X"00",
56543=>X"00",
56544=>X"00",
56545=>X"00",
56546=>X"00",
56547=>X"00",
56548=>X"00",
56549=>X"00",
56550=>X"00",
56551=>X"00",
56552=>X"00",
56553=>X"00",
56554=>X"00",
56555=>X"00",
56556=>X"00",
56557=>X"00",
56558=>X"00",
56559=>X"00",
56560=>X"00",
56561=>X"00",
56562=>X"00",
56563=>X"00",
56564=>X"00",
56565=>X"00",
56566=>X"00",
56567=>X"00",
56568=>X"00",
56569=>X"00",
56570=>X"00",
56571=>X"00",
56572=>X"00",
56573=>X"00",
56574=>X"00",
56575=>X"00",
56576=>X"00",
56577=>X"00",
56578=>X"00",
56579=>X"00",
56580=>X"00",
56581=>X"00",
56582=>X"00",
56583=>X"00",
56584=>X"00",
56585=>X"00",
56586=>X"00",
56587=>X"00",
56588=>X"00",
56589=>X"00",
56590=>X"00",
56591=>X"00",
56592=>X"00",
56593=>X"00",
56594=>X"00",
56595=>X"00",
56596=>X"00",
56597=>X"00",
56598=>X"00",
56599=>X"00",
56600=>X"00",
56601=>X"00",
56602=>X"00",
56603=>X"00",
56604=>X"00",
56605=>X"00",
56606=>X"00",
56607=>X"00",
56608=>X"00",
56609=>X"00",
56610=>X"00",
56611=>X"00",
56612=>X"00",
56613=>X"00",
56614=>X"00",
56615=>X"00",
56616=>X"00",
56617=>X"00",
56618=>X"00",
56619=>X"00",
56620=>X"00",
56621=>X"00",
56622=>X"00",
56623=>X"00",
56624=>X"00",
56625=>X"00",
56626=>X"00",
56627=>X"00",
56628=>X"00",
56629=>X"00",
56630=>X"00",
56631=>X"00",
56632=>X"00",
56633=>X"00",
56634=>X"00",
56635=>X"00",
56636=>X"00",
56637=>X"00",
56638=>X"00",
56639=>X"00",
56640=>X"00",
56641=>X"00",
56642=>X"00",
56643=>X"00",
56644=>X"00",
56645=>X"00",
56646=>X"00",
56647=>X"00",
56648=>X"00",
56649=>X"00",
56650=>X"00",
56651=>X"00",
56652=>X"00",
56653=>X"00",
56654=>X"00",
56655=>X"00",
56656=>X"00",
56657=>X"00",
56658=>X"00",
56659=>X"00",
56660=>X"00",
56661=>X"00",
56662=>X"00",
56663=>X"00",
56664=>X"00",
56665=>X"00",
56666=>X"00",
56667=>X"00",
56668=>X"00",
56669=>X"00",
56670=>X"00",
56671=>X"00",
56672=>X"00",
56673=>X"00",
56674=>X"00",
56675=>X"00",
56676=>X"00",
56677=>X"00",
56678=>X"00",
56679=>X"00",
56680=>X"00",
56681=>X"00",
56682=>X"00",
56683=>X"00",
56684=>X"00",
56685=>X"00",
56686=>X"00",
56687=>X"00",
56688=>X"00",
56689=>X"00",
56690=>X"00",
56691=>X"00",
56692=>X"00",
56693=>X"00",
56694=>X"00",
56695=>X"00",
56696=>X"00",
56697=>X"00",
56698=>X"00",
56699=>X"00",
56700=>X"00",
56701=>X"00",
56702=>X"00",
56703=>X"00",
56704=>X"00",
56705=>X"00",
56706=>X"00",
56707=>X"00",
56708=>X"00",
56709=>X"00",
56710=>X"00",
56711=>X"00",
56712=>X"00",
56713=>X"00",
56714=>X"00",
56715=>X"00",
56716=>X"00",
56717=>X"00",
56718=>X"00",
56719=>X"00",
56720=>X"00",
56721=>X"00",
56722=>X"00",
56723=>X"00",
56724=>X"00",
56725=>X"00",
56726=>X"00",
56727=>X"00",
56728=>X"00",
56729=>X"00",
56730=>X"00",
56731=>X"00",
56732=>X"00",
56733=>X"00",
56734=>X"00",
56735=>X"00",
56736=>X"00",
56737=>X"00",
56738=>X"00",
56739=>X"00",
56740=>X"00",
56741=>X"00",
56742=>X"00",
56743=>X"00",
56744=>X"00",
56745=>X"00",
56746=>X"00",
56747=>X"00",
56748=>X"00",
56749=>X"00",
56750=>X"00",
56751=>X"00",
56752=>X"00",
56753=>X"00",
56754=>X"00",
56755=>X"00",
56756=>X"00",
56757=>X"00",
56758=>X"00",
56759=>X"00",
56760=>X"00",
56761=>X"00",
56762=>X"00",
56763=>X"00",
56764=>X"00",
56765=>X"00",
56766=>X"00",
56767=>X"00",
56768=>X"00",
56769=>X"00",
56770=>X"00",
56771=>X"00",
56772=>X"00",
56773=>X"00",
56774=>X"00",
56775=>X"00",
56776=>X"00",
56777=>X"00",
56778=>X"00",
56779=>X"00",
56780=>X"00",
56781=>X"00",
56782=>X"00",
56783=>X"00",
56784=>X"00",
56785=>X"00",
56786=>X"00",
56787=>X"00",
56788=>X"00",
56789=>X"00",
56790=>X"00",
56791=>X"00",
56792=>X"00",
56793=>X"00",
56794=>X"00",
56795=>X"00",
56796=>X"00",
56797=>X"00",
56798=>X"00",
56799=>X"00",
56800=>X"00",
56801=>X"00",
56802=>X"00",
56803=>X"00",
56804=>X"00",
56805=>X"00",
56806=>X"00",
56807=>X"00",
56808=>X"00",
56809=>X"00",
56810=>X"00",
56811=>X"00",
56812=>X"00",
56813=>X"00",
56814=>X"00",
56815=>X"00",
56816=>X"00",
56817=>X"00",
56818=>X"00",
56819=>X"00",
56820=>X"00",
56821=>X"00",
56822=>X"00",
56823=>X"00",
56824=>X"00",
56825=>X"00",
56826=>X"00",
56827=>X"00",
56828=>X"00",
56829=>X"00",
56830=>X"00",
56831=>X"00",
56832=>X"00",
56833=>X"00",
56834=>X"00",
56835=>X"00",
56836=>X"00",
56837=>X"00",
56838=>X"00",
56839=>X"00",
56840=>X"00",
56841=>X"00",
56842=>X"00",
56843=>X"00",
56844=>X"00",
56845=>X"00",
56846=>X"00",
56847=>X"00",
56848=>X"00",
56849=>X"00",
56850=>X"00",
56851=>X"00",
56852=>X"00",
56853=>X"00",
56854=>X"00",
56855=>X"00",
56856=>X"00",
56857=>X"00",
56858=>X"00",
56859=>X"00",
56860=>X"00",
56861=>X"00",
56862=>X"00",
56863=>X"00",
56864=>X"00",
56865=>X"00",
56866=>X"00",
56867=>X"00",
56868=>X"00",
56869=>X"00",
56870=>X"00",
56871=>X"00",
56872=>X"00",
56873=>X"00",
56874=>X"00",
56875=>X"00",
56876=>X"00",
56877=>X"00",
56878=>X"00",
56879=>X"00",
56880=>X"00",
56881=>X"00",
56882=>X"00",
56883=>X"00",
56884=>X"00",
56885=>X"00",
56886=>X"00",
56887=>X"00",
56888=>X"00",
56889=>X"00",
56890=>X"00",
56891=>X"00",
56892=>X"00",
56893=>X"00",
56894=>X"00",
56895=>X"00",
56896=>X"00",
56897=>X"00",
56898=>X"00",
56899=>X"00",
56900=>X"00",
56901=>X"00",
56902=>X"00",
56903=>X"00",
56904=>X"00",
56905=>X"00",
56906=>X"00",
56907=>X"00",
56908=>X"00",
56909=>X"00",
56910=>X"00",
56911=>X"00",
56912=>X"00",
56913=>X"00",
56914=>X"00",
56915=>X"00",
56916=>X"00",
56917=>X"00",
56918=>X"00",
56919=>X"00",
56920=>X"00",
56921=>X"00",
56922=>X"00",
56923=>X"00",
56924=>X"00",
56925=>X"00",
56926=>X"00",
56927=>X"00",
56928=>X"00",
56929=>X"00",
56930=>X"00",
56931=>X"00",
56932=>X"00",
56933=>X"00",
56934=>X"00",
56935=>X"00",
56936=>X"00",
56937=>X"00",
56938=>X"00",
56939=>X"00",
56940=>X"00",
56941=>X"00",
56942=>X"00",
56943=>X"00",
56944=>X"00",
56945=>X"00",
56946=>X"00",
56947=>X"00",
56948=>X"00",
56949=>X"00",
56950=>X"00",
56951=>X"00",
56952=>X"00",
56953=>X"00",
56954=>X"00",
56955=>X"00",
56956=>X"00",
56957=>X"00",
56958=>X"00",
56959=>X"00",
56960=>X"00",
56961=>X"00",
56962=>X"00",
56963=>X"00",
56964=>X"00",
56965=>X"00",
56966=>X"00",
56967=>X"00",
56968=>X"00",
56969=>X"00",
56970=>X"00",
56971=>X"00",
56972=>X"00",
56973=>X"00",
56974=>X"00",
56975=>X"00",
56976=>X"00",
56977=>X"00",
56978=>X"00",
56979=>X"00",
56980=>X"00",
56981=>X"00",
56982=>X"00",
56983=>X"00",
56984=>X"00",
56985=>X"00",
56986=>X"00",
56987=>X"00",
56988=>X"00",
56989=>X"00",
56990=>X"00",
56991=>X"00",
56992=>X"00",
56993=>X"00",
56994=>X"00",
56995=>X"00",
56996=>X"00",
56997=>X"00",
56998=>X"00",
56999=>X"00",
57000=>X"00",
57001=>X"00",
57002=>X"00",
57003=>X"00",
57004=>X"00",
57005=>X"00",
57006=>X"00",
57007=>X"00",
57008=>X"00",
57009=>X"00",
57010=>X"00",
57011=>X"00",
57012=>X"00",
57013=>X"00",
57014=>X"00",
57015=>X"00",
57016=>X"00",
57017=>X"00",
57018=>X"00",
57019=>X"00",
57020=>X"00",
57021=>X"00",
57022=>X"00",
57023=>X"00",
57024=>X"00",
57025=>X"00",
57026=>X"00",
57027=>X"00",
57028=>X"00",
57029=>X"00",
57030=>X"00",
57031=>X"00",
57032=>X"00",
57033=>X"00",
57034=>X"00",
57035=>X"00",
57036=>X"00",
57037=>X"00",
57038=>X"00",
57039=>X"00",
57040=>X"00",
57041=>X"00",
57042=>X"00",
57043=>X"00",
57044=>X"00",
57045=>X"00",
57046=>X"00",
57047=>X"00",
57048=>X"00",
57049=>X"00",
57050=>X"00",
57051=>X"00",
57052=>X"00",
57053=>X"00",
57054=>X"00",
57055=>X"00",
57056=>X"00",
57057=>X"00",
57058=>X"00",
57059=>X"00",
57060=>X"00",
57061=>X"00",
57062=>X"00",
57063=>X"00",
57064=>X"00",
57065=>X"00",
57066=>X"00",
57067=>X"00",
57068=>X"00",
57069=>X"00",
57070=>X"00",
57071=>X"00",
57072=>X"00",
57073=>X"00",
57074=>X"00",
57075=>X"00",
57076=>X"00",
57077=>X"00",
57078=>X"00",
57079=>X"00",
57080=>X"00",
57081=>X"00",
57082=>X"00",
57083=>X"00",
57084=>X"00",
57085=>X"00",
57086=>X"00",
57087=>X"00",
57088=>X"00",
57089=>X"00",
57090=>X"00",
57091=>X"00",
57092=>X"00",
57093=>X"00",
57094=>X"00",
57095=>X"00",
57096=>X"00",
57097=>X"00",
57098=>X"00",
57099=>X"00",
57100=>X"00",
57101=>X"00",
57102=>X"00",
57103=>X"00",
57104=>X"00",
57105=>X"00",
57106=>X"00",
57107=>X"00",
57108=>X"00",
57109=>X"00",
57110=>X"00",
57111=>X"00",
57112=>X"00",
57113=>X"00",
57114=>X"00",
57115=>X"00",
57116=>X"00",
57117=>X"00",
57118=>X"00",
57119=>X"00",
57120=>X"00",
57121=>X"00",
57122=>X"00",
57123=>X"00",
57124=>X"00",
57125=>X"00",
57126=>X"00",
57127=>X"00",
57128=>X"00",
57129=>X"00",
57130=>X"00",
57131=>X"00",
57132=>X"00",
57133=>X"00",
57134=>X"00",
57135=>X"00",
57136=>X"00",
57137=>X"00",
57138=>X"00",
57139=>X"00",
57140=>X"00",
57141=>X"00",
57142=>X"00",
57143=>X"00",
57144=>X"00",
57145=>X"00",
57146=>X"00",
57147=>X"00",
57148=>X"00",
57149=>X"00",
57150=>X"00",
57151=>X"00",
57152=>X"00",
57153=>X"00",
57154=>X"00",
57155=>X"00",
57156=>X"00",
57157=>X"00",
57158=>X"00",
57159=>X"00",
57160=>X"00",
57161=>X"00",
57162=>X"00",
57163=>X"00",
57164=>X"00",
57165=>X"00",
57166=>X"00",
57167=>X"00",
57168=>X"00",
57169=>X"00",
57170=>X"00",
57171=>X"00",
57172=>X"00",
57173=>X"00",
57174=>X"00",
57175=>X"00",
57176=>X"00",
57177=>X"00",
57178=>X"00",
57179=>X"00",
57180=>X"00",
57181=>X"00",
57182=>X"00",
57183=>X"00",
57184=>X"00",
57185=>X"00",
57186=>X"00",
57187=>X"00",
57188=>X"00",
57189=>X"00",
57190=>X"00",
57191=>X"00",
57192=>X"00",
57193=>X"00",
57194=>X"00",
57195=>X"00",
57196=>X"00",
57197=>X"00",
57198=>X"00",
57199=>X"00",
57200=>X"00",
57201=>X"00",
57202=>X"00",
57203=>X"00",
57204=>X"00",
57205=>X"00",
57206=>X"00",
57207=>X"00",
57208=>X"00",
57209=>X"00",
57210=>X"00",
57211=>X"00",
57212=>X"00",
57213=>X"00",
57214=>X"00",
57215=>X"00",
57216=>X"00",
57217=>X"00",
57218=>X"00",
57219=>X"00",
57220=>X"00",
57221=>X"00",
57222=>X"00",
57223=>X"00",
57224=>X"00",
57225=>X"00",
57226=>X"00",
57227=>X"00",
57228=>X"00",
57229=>X"00",
57230=>X"00",
57231=>X"00",
57232=>X"00",
57233=>X"00",
57234=>X"00",
57235=>X"00",
57236=>X"00",
57237=>X"00",
57238=>X"00",
57239=>X"00",
57240=>X"00",
57241=>X"00",
57242=>X"00",
57243=>X"00",
57244=>X"00",
57245=>X"00",
57246=>X"00",
57247=>X"00",
57248=>X"00",
57249=>X"00",
57250=>X"00",
57251=>X"00",
57252=>X"00",
57253=>X"00",
57254=>X"00",
57255=>X"00",
57256=>X"00",
57257=>X"00",
57258=>X"00",
57259=>X"00",
57260=>X"00",
57261=>X"00",
57262=>X"00",
57263=>X"00",
57264=>X"00",
57265=>X"00",
57266=>X"00",
57267=>X"00",
57268=>X"00",
57269=>X"00",
57270=>X"00",
57271=>X"00",
57272=>X"00",
57273=>X"00",
57274=>X"00",
57275=>X"00",
57276=>X"00",
57277=>X"00",
57278=>X"00",
57279=>X"00",
57280=>X"00",
57281=>X"00",
57282=>X"00",
57283=>X"00",
57284=>X"00",
57285=>X"00",
57286=>X"00",
57287=>X"00",
57288=>X"00",
57289=>X"00",
57290=>X"00",
57291=>X"00",
57292=>X"00",
57293=>X"00",
57294=>X"00",
57295=>X"00",
57296=>X"00",
57297=>X"00",
57298=>X"00",
57299=>X"00",
57300=>X"00",
57301=>X"00",
57302=>X"00",
57303=>X"00",
57304=>X"00",
57305=>X"00",
57306=>X"00",
57307=>X"00",
57308=>X"00",
57309=>X"00",
57310=>X"00",
57311=>X"00",
57312=>X"00",
57313=>X"00",
57314=>X"00",
57315=>X"00",
57316=>X"00",
57317=>X"00",
57318=>X"00",
57319=>X"00",
57320=>X"00",
57321=>X"00",
57322=>X"00",
57323=>X"00",
57324=>X"00",
57325=>X"00",
57326=>X"00",
57327=>X"00",
57328=>X"00",
57329=>X"00",
57330=>X"00",
57331=>X"00",
57332=>X"00",
57333=>X"00",
57334=>X"00",
57335=>X"00",
57336=>X"00",
57337=>X"00",
57338=>X"00",
57339=>X"00",
57340=>X"00",
57341=>X"00",
57342=>X"00",
57343=>X"00",
57344=>X"00",
57345=>X"00",
57346=>X"00",
57347=>X"00",
57348=>X"00",
57349=>X"00",
57350=>X"00",
57351=>X"00",
57352=>X"00",
57353=>X"00",
57354=>X"00",
57355=>X"00",
57356=>X"00",
57357=>X"00",
57358=>X"00",
57359=>X"00",
57360=>X"00",
57361=>X"00",
57362=>X"00",
57363=>X"00",
57364=>X"00",
57365=>X"00",
57366=>X"00",
57367=>X"00",
57368=>X"00",
57369=>X"00",
57370=>X"00",
57371=>X"00",
57372=>X"00",
57373=>X"00",
57374=>X"00",
57375=>X"00",
57376=>X"00",
57377=>X"00",
57378=>X"00",
57379=>X"00",
57380=>X"00",
57381=>X"00",
57382=>X"00",
57383=>X"00",
57384=>X"00",
57385=>X"00",
57386=>X"00",
57387=>X"00",
57388=>X"00",
57389=>X"00",
57390=>X"00",
57391=>X"00",
57392=>X"00",
57393=>X"00",
57394=>X"00",
57395=>X"00",
57396=>X"00",
57397=>X"00",
57398=>X"00",
57399=>X"00",
57400=>X"00",
57401=>X"00",
57402=>X"00",
57403=>X"00",
57404=>X"00",
57405=>X"00",
57406=>X"00",
57407=>X"00",
57408=>X"00",
57409=>X"00",
57410=>X"00",
57411=>X"00",
57412=>X"00",
57413=>X"00",
57414=>X"00",
57415=>X"00",
57416=>X"00",
57417=>X"00",
57418=>X"00",
57419=>X"00",
57420=>X"00",
57421=>X"00",
57422=>X"00",
57423=>X"00",
57424=>X"00",
57425=>X"00",
57426=>X"00",
57427=>X"00",
57428=>X"00",
57429=>X"00",
57430=>X"00",
57431=>X"00",
57432=>X"00",
57433=>X"00",
57434=>X"00",
57435=>X"00",
57436=>X"00",
57437=>X"00",
57438=>X"00",
57439=>X"00",
57440=>X"00",
57441=>X"00",
57442=>X"00",
57443=>X"00",
57444=>X"00",
57445=>X"00",
57446=>X"00",
57447=>X"00",
57448=>X"00",
57449=>X"00",
57450=>X"00",
57451=>X"00",
57452=>X"00",
57453=>X"00",
57454=>X"00",
57455=>X"00",
57456=>X"00",
57457=>X"00",
57458=>X"00",
57459=>X"00",
57460=>X"00",
57461=>X"00",
57462=>X"00",
57463=>X"00",
57464=>X"00",
57465=>X"00",
57466=>X"00",
57467=>X"00",
57468=>X"00",
57469=>X"00",
57470=>X"00",
57471=>X"00",
57472=>X"00",
57473=>X"00",
57474=>X"00",
57475=>X"00",
57476=>X"00",
57477=>X"00",
57478=>X"00",
57479=>X"00",
57480=>X"00",
57481=>X"00",
57482=>X"00",
57483=>X"00",
57484=>X"00",
57485=>X"00",
57486=>X"00",
57487=>X"00",
57488=>X"00",
57489=>X"00",
57490=>X"00",
57491=>X"00",
57492=>X"00",
57493=>X"00",
57494=>X"00",
57495=>X"00",
57496=>X"00",
57497=>X"00",
57498=>X"00",
57499=>X"00",
57500=>X"00",
57501=>X"00",
57502=>X"00",
57503=>X"00",
57504=>X"00",
57505=>X"00",
57506=>X"00",
57507=>X"00",
57508=>X"00",
57509=>X"00",
57510=>X"00",
57511=>X"00",
57512=>X"00",
57513=>X"00",
57514=>X"00",
57515=>X"00",
57516=>X"00",
57517=>X"00",
57518=>X"00",
57519=>X"00",
57520=>X"00",
57521=>X"00",
57522=>X"00",
57523=>X"00",
57524=>X"00",
57525=>X"00",
57526=>X"00",
57527=>X"00",
57528=>X"00",
57529=>X"00",
57530=>X"00",
57531=>X"00",
57532=>X"00",
57533=>X"00",
57534=>X"00",
57535=>X"00",
57536=>X"00",
57537=>X"00",
57538=>X"00",
57539=>X"00",
57540=>X"00",
57541=>X"00",
57542=>X"00",
57543=>X"00",
57544=>X"00",
57545=>X"00",
57546=>X"00",
57547=>X"00",
57548=>X"00",
57549=>X"00",
57550=>X"00",
57551=>X"00",
57552=>X"00",
57553=>X"00",
57554=>X"00",
57555=>X"00",
57556=>X"00",
57557=>X"00",
57558=>X"00",
57559=>X"00",
57560=>X"00",
57561=>X"00",
57562=>X"00",
57563=>X"00",
57564=>X"00",
57565=>X"00",
57566=>X"00",
57567=>X"00",
57568=>X"00",
57569=>X"00",
57570=>X"00",
57571=>X"00",
57572=>X"00",
57573=>X"00",
57574=>X"00",
57575=>X"00",
57576=>X"00",
57577=>X"00",
57578=>X"00",
57579=>X"00",
57580=>X"00",
57581=>X"00",
57582=>X"00",
57583=>X"00",
57584=>X"00",
57585=>X"00",
57586=>X"00",
57587=>X"00",
57588=>X"00",
57589=>X"00",
57590=>X"00",
57591=>X"00",
57592=>X"00",
57593=>X"00",
57594=>X"00",
57595=>X"00",
57596=>X"00",
57597=>X"00",
57598=>X"00",
57599=>X"00",
57600=>X"00",
57601=>X"00",
57602=>X"00",
57603=>X"00",
57604=>X"00",
57605=>X"00",
57606=>X"00",
57607=>X"00",
57608=>X"00",
57609=>X"00",
57610=>X"00",
57611=>X"00",
57612=>X"00",
57613=>X"00",
57614=>X"00",
57615=>X"00",
57616=>X"00",
57617=>X"00",
57618=>X"00",
57619=>X"00",
57620=>X"00",
57621=>X"00",
57622=>X"00",
57623=>X"00",
57624=>X"00",
57625=>X"00",
57626=>X"00",
57627=>X"00",
57628=>X"00",
57629=>X"00",
57630=>X"00",
57631=>X"00",
57632=>X"00",
57633=>X"00",
57634=>X"00",
57635=>X"00",
57636=>X"00",
57637=>X"00",
57638=>X"00",
57639=>X"00",
57640=>X"00",
57641=>X"00",
57642=>X"00",
57643=>X"00",
57644=>X"00",
57645=>X"00",
57646=>X"00",
57647=>X"00",
57648=>X"00",
57649=>X"00",
57650=>X"00",
57651=>X"00",
57652=>X"00",
57653=>X"00",
57654=>X"00",
57655=>X"00",
57656=>X"00",
57657=>X"00",
57658=>X"00",
57659=>X"00",
57660=>X"00",
57661=>X"00",
57662=>X"00",
57663=>X"00",
57664=>X"00",
57665=>X"00",
57666=>X"00",
57667=>X"00",
57668=>X"00",
57669=>X"00",
57670=>X"00",
57671=>X"00",
57672=>X"00",
57673=>X"00",
57674=>X"00",
57675=>X"00",
57676=>X"00",
57677=>X"00",
57678=>X"00",
57679=>X"00",
57680=>X"00",
57681=>X"00",
57682=>X"00",
57683=>X"00",
57684=>X"00",
57685=>X"00",
57686=>X"00",
57687=>X"00",
57688=>X"00",
57689=>X"00",
57690=>X"00",
57691=>X"00",
57692=>X"00",
57693=>X"00",
57694=>X"00",
57695=>X"00",
57696=>X"00",
57697=>X"00",
57698=>X"00",
57699=>X"00",
57700=>X"00",
57701=>X"00",
57702=>X"00",
57703=>X"00",
57704=>X"00",
57705=>X"00",
57706=>X"00",
57707=>X"00",
57708=>X"00",
57709=>X"00",
57710=>X"00",
57711=>X"00",
57712=>X"00",
57713=>X"00",
57714=>X"00",
57715=>X"00",
57716=>X"00",
57717=>X"00",
57718=>X"00",
57719=>X"00",
57720=>X"00",
57721=>X"00",
57722=>X"00",
57723=>X"00",
57724=>X"00",
57725=>X"00",
57726=>X"00",
57727=>X"00",
57728=>X"00",
57729=>X"00",
57730=>X"00",
57731=>X"00",
57732=>X"00",
57733=>X"00",
57734=>X"00",
57735=>X"00",
57736=>X"00",
57737=>X"00",
57738=>X"00",
57739=>X"00",
57740=>X"00",
57741=>X"00",
57742=>X"00",
57743=>X"00",
57744=>X"00",
57745=>X"00",
57746=>X"00",
57747=>X"00",
57748=>X"00",
57749=>X"00",
57750=>X"00",
57751=>X"00",
57752=>X"00",
57753=>X"00",
57754=>X"00",
57755=>X"00",
57756=>X"00",
57757=>X"00",
57758=>X"00",
57759=>X"00",
57760=>X"00",
57761=>X"00",
57762=>X"00",
57763=>X"00",
57764=>X"00",
57765=>X"00",
57766=>X"00",
57767=>X"00",
57768=>X"00",
57769=>X"00",
57770=>X"00",
57771=>X"00",
57772=>X"00",
57773=>X"00",
57774=>X"00",
57775=>X"00",
57776=>X"00",
57777=>X"00",
57778=>X"00",
57779=>X"00",
57780=>X"00",
57781=>X"00",
57782=>X"00",
57783=>X"00",
57784=>X"00",
57785=>X"00",
57786=>X"00",
57787=>X"00",
57788=>X"00",
57789=>X"00",
57790=>X"00",
57791=>X"00",
57792=>X"00",
57793=>X"00",
57794=>X"00",
57795=>X"00",
57796=>X"00",
57797=>X"00",
57798=>X"00",
57799=>X"00",
57800=>X"00",
57801=>X"00",
57802=>X"00",
57803=>X"00",
57804=>X"00",
57805=>X"00",
57806=>X"00",
57807=>X"00",
57808=>X"00",
57809=>X"00",
57810=>X"00",
57811=>X"00",
57812=>X"00",
57813=>X"00",
57814=>X"00",
57815=>X"00",
57816=>X"00",
57817=>X"00",
57818=>X"00",
57819=>X"00",
57820=>X"00",
57821=>X"00",
57822=>X"00",
57823=>X"00",
57824=>X"00",
57825=>X"00",
57826=>X"00",
57827=>X"00",
57828=>X"00",
57829=>X"00",
57830=>X"00",
57831=>X"00",
57832=>X"00",
57833=>X"00",
57834=>X"00",
57835=>X"00",
57836=>X"00",
57837=>X"00",
57838=>X"00",
57839=>X"00",
57840=>X"00",
57841=>X"00",
57842=>X"00",
57843=>X"00",
57844=>X"00",
57845=>X"00",
57846=>X"00",
57847=>X"00",
57848=>X"00",
57849=>X"00",
57850=>X"00",
57851=>X"00",
57852=>X"00",
57853=>X"00",
57854=>X"00",
57855=>X"00",
57856=>X"00",
57857=>X"00",
57858=>X"00",
57859=>X"00",
57860=>X"00",
57861=>X"00",
57862=>X"00",
57863=>X"00",
57864=>X"00",
57865=>X"00",
57866=>X"00",
57867=>X"00",
57868=>X"00",
57869=>X"00",
57870=>X"00",
57871=>X"00",
57872=>X"00",
57873=>X"00",
57874=>X"00",
57875=>X"00",
57876=>X"00",
57877=>X"00",
57878=>X"00",
57879=>X"00",
57880=>X"00",
57881=>X"00",
57882=>X"00",
57883=>X"00",
57884=>X"00",
57885=>X"00",
57886=>X"00",
57887=>X"00",
57888=>X"00",
57889=>X"00",
57890=>X"00",
57891=>X"00",
57892=>X"00",
57893=>X"00",
57894=>X"00",
57895=>X"00",
57896=>X"00",
57897=>X"00",
57898=>X"00",
57899=>X"00",
57900=>X"00",
57901=>X"00",
57902=>X"00",
57903=>X"00",
57904=>X"00",
57905=>X"00",
57906=>X"00",
57907=>X"00",
57908=>X"00",
57909=>X"00",
57910=>X"00",
57911=>X"00",
57912=>X"00",
57913=>X"00",
57914=>X"00",
57915=>X"00",
57916=>X"00",
57917=>X"00",
57918=>X"00",
57919=>X"00",
57920=>X"00",
57921=>X"00",
57922=>X"00",
57923=>X"00",
57924=>X"00",
57925=>X"00",
57926=>X"00",
57927=>X"00",
57928=>X"00",
57929=>X"00",
57930=>X"00",
57931=>X"00",
57932=>X"00",
57933=>X"00",
57934=>X"00",
57935=>X"00",
57936=>X"00",
57937=>X"00",
57938=>X"00",
57939=>X"00",
57940=>X"00",
57941=>X"00",
57942=>X"00",
57943=>X"00",
57944=>X"00",
57945=>X"00",
57946=>X"00",
57947=>X"00",
57948=>X"00",
57949=>X"00",
57950=>X"00",
57951=>X"00",
57952=>X"00",
57953=>X"00",
57954=>X"00",
57955=>X"00",
57956=>X"00",
57957=>X"00",
57958=>X"00",
57959=>X"00",
57960=>X"00",
57961=>X"00",
57962=>X"00",
57963=>X"00",
57964=>X"00",
57965=>X"00",
57966=>X"00",
57967=>X"00",
57968=>X"00",
57969=>X"00",
57970=>X"00",
57971=>X"00",
57972=>X"00",
57973=>X"00",
57974=>X"00",
57975=>X"00",
57976=>X"00",
57977=>X"00",
57978=>X"00",
57979=>X"00",
57980=>X"00",
57981=>X"00",
57982=>X"00",
57983=>X"00",
57984=>X"00",
57985=>X"00",
57986=>X"00",
57987=>X"00",
57988=>X"00",
57989=>X"00",
57990=>X"00",
57991=>X"00",
57992=>X"00",
57993=>X"00",
57994=>X"00",
57995=>X"00",
57996=>X"00",
57997=>X"00",
57998=>X"00",
57999=>X"00",
58000=>X"00",
58001=>X"00",
58002=>X"00",
58003=>X"00",
58004=>X"00",
58005=>X"00",
58006=>X"00",
58007=>X"00",
58008=>X"00",
58009=>X"00",
58010=>X"00",
58011=>X"00",
58012=>X"00",
58013=>X"00",
58014=>X"00",
58015=>X"00",
58016=>X"00",
58017=>X"00",
58018=>X"00",
58019=>X"00",
58020=>X"00",
58021=>X"00",
58022=>X"00",
58023=>X"00",
58024=>X"00",
58025=>X"00",
58026=>X"00",
58027=>X"00",
58028=>X"00",
58029=>X"00",
58030=>X"00",
58031=>X"00",
58032=>X"00",
58033=>X"00",
58034=>X"00",
58035=>X"00",
58036=>X"00",
58037=>X"00",
58038=>X"00",
58039=>X"00",
58040=>X"00",
58041=>X"00",
58042=>X"00",
58043=>X"00",
58044=>X"00",
58045=>X"00",
58046=>X"00",
58047=>X"00",
58048=>X"00",
58049=>X"00",
58050=>X"00",
58051=>X"00",
58052=>X"00",
58053=>X"00",
58054=>X"00",
58055=>X"00",
58056=>X"00",
58057=>X"00",
58058=>X"00",
58059=>X"00",
58060=>X"00",
58061=>X"00",
58062=>X"00",
58063=>X"00",
58064=>X"00",
58065=>X"00",
58066=>X"00",
58067=>X"00",
58068=>X"00",
58069=>X"00",
58070=>X"00",
58071=>X"00",
58072=>X"00",
58073=>X"00",
58074=>X"00",
58075=>X"00",
58076=>X"00",
58077=>X"00",
58078=>X"00",
58079=>X"00",
58080=>X"00",
58081=>X"00",
58082=>X"00",
58083=>X"00",
58084=>X"00",
58085=>X"00",
58086=>X"00",
58087=>X"00",
58088=>X"00",
58089=>X"00",
58090=>X"00",
58091=>X"00",
58092=>X"00",
58093=>X"00",
58094=>X"00",
58095=>X"00",
58096=>X"00",
58097=>X"00",
58098=>X"00",
58099=>X"00",
58100=>X"00",
58101=>X"00",
58102=>X"00",
58103=>X"00",
58104=>X"00",
58105=>X"00",
58106=>X"00",
58107=>X"00",
58108=>X"00",
58109=>X"00",
58110=>X"00",
58111=>X"00",
58112=>X"00",
58113=>X"00",
58114=>X"00",
58115=>X"00",
58116=>X"00",
58117=>X"00",
58118=>X"00",
58119=>X"00",
58120=>X"00",
58121=>X"00",
58122=>X"00",
58123=>X"00",
58124=>X"00",
58125=>X"00",
58126=>X"00",
58127=>X"00",
58128=>X"00",
58129=>X"00",
58130=>X"00",
58131=>X"00",
58132=>X"00",
58133=>X"00",
58134=>X"00",
58135=>X"00",
58136=>X"00",
58137=>X"00",
58138=>X"00",
58139=>X"00",
58140=>X"00",
58141=>X"00",
58142=>X"00",
58143=>X"00",
58144=>X"00",
58145=>X"00",
58146=>X"00",
58147=>X"00",
58148=>X"00",
58149=>X"00",
58150=>X"00",
58151=>X"00",
58152=>X"00",
58153=>X"00",
58154=>X"00",
58155=>X"00",
58156=>X"00",
58157=>X"00",
58158=>X"00",
58159=>X"00",
58160=>X"00",
58161=>X"00",
58162=>X"00",
58163=>X"00",
58164=>X"00",
58165=>X"00",
58166=>X"00",
58167=>X"00",
58168=>X"00",
58169=>X"00",
58170=>X"00",
58171=>X"00",
58172=>X"00",
58173=>X"00",
58174=>X"00",
58175=>X"00",
58176=>X"00",
58177=>X"00",
58178=>X"00",
58179=>X"00",
58180=>X"00",
58181=>X"00",
58182=>X"00",
58183=>X"00",
58184=>X"00",
58185=>X"00",
58186=>X"00",
58187=>X"00",
58188=>X"00",
58189=>X"00",
58190=>X"00",
58191=>X"00",
58192=>X"00",
58193=>X"00",
58194=>X"00",
58195=>X"00",
58196=>X"00",
58197=>X"00",
58198=>X"00",
58199=>X"00",
58200=>X"00",
58201=>X"00",
58202=>X"00",
58203=>X"00",
58204=>X"00",
58205=>X"00",
58206=>X"00",
58207=>X"00",
58208=>X"00",
58209=>X"00",
58210=>X"00",
58211=>X"00",
58212=>X"00",
58213=>X"00",
58214=>X"00",
58215=>X"00",
58216=>X"00",
58217=>X"00",
58218=>X"00",
58219=>X"00",
58220=>X"00",
58221=>X"00",
58222=>X"00",
58223=>X"00",
58224=>X"00",
58225=>X"00",
58226=>X"00",
58227=>X"00",
58228=>X"00",
58229=>X"00",
58230=>X"00",
58231=>X"00",
58232=>X"00",
58233=>X"00",
58234=>X"00",
58235=>X"00",
58236=>X"00",
58237=>X"00",
58238=>X"00",
58239=>X"00",
58240=>X"00",
58241=>X"00",
58242=>X"00",
58243=>X"00",
58244=>X"00",
58245=>X"00",
58246=>X"00",
58247=>X"00",
58248=>X"00",
58249=>X"00",
58250=>X"00",
58251=>X"00",
58252=>X"00",
58253=>X"00",
58254=>X"00",
58255=>X"00",
58256=>X"00",
58257=>X"00",
58258=>X"00",
58259=>X"00",
58260=>X"00",
58261=>X"00",
58262=>X"00",
58263=>X"00",
58264=>X"00",
58265=>X"00",
58266=>X"00",
58267=>X"00",
58268=>X"00",
58269=>X"00",
58270=>X"00",
58271=>X"00",
58272=>X"00",
58273=>X"00",
58274=>X"00",
58275=>X"00",
58276=>X"00",
58277=>X"00",
58278=>X"00",
58279=>X"00",
58280=>X"00",
58281=>X"00",
58282=>X"00",
58283=>X"00",
58284=>X"00",
58285=>X"00",
58286=>X"00",
58287=>X"00",
58288=>X"00",
58289=>X"00",
58290=>X"00",
58291=>X"00",
58292=>X"00",
58293=>X"00",
58294=>X"00",
58295=>X"00",
58296=>X"00",
58297=>X"00",
58298=>X"00",
58299=>X"00",
58300=>X"00",
58301=>X"00",
58302=>X"00",
58303=>X"00",
58304=>X"00",
58305=>X"00",
58306=>X"00",
58307=>X"00",
58308=>X"00",
58309=>X"00",
58310=>X"00",
58311=>X"00",
58312=>X"00",
58313=>X"00",
58314=>X"00",
58315=>X"00",
58316=>X"00",
58317=>X"00",
58318=>X"00",
58319=>X"00",
58320=>X"00",
58321=>X"00",
58322=>X"00",
58323=>X"00",
58324=>X"00",
58325=>X"00",
58326=>X"00",
58327=>X"00",
58328=>X"00",
58329=>X"00",
58330=>X"00",
58331=>X"00",
58332=>X"00",
58333=>X"00",
58334=>X"00",
58335=>X"00",
58336=>X"00",
58337=>X"00",
58338=>X"00",
58339=>X"00",
58340=>X"00",
58341=>X"00",
58342=>X"00",
58343=>X"00",
58344=>X"00",
58345=>X"00",
58346=>X"00",
58347=>X"00",
58348=>X"00",
58349=>X"00",
58350=>X"00",
58351=>X"00",
58352=>X"00",
58353=>X"00",
58354=>X"00",
58355=>X"00",
58356=>X"00",
58357=>X"00",
58358=>X"00",
58359=>X"00",
58360=>X"00",
58361=>X"00",
58362=>X"00",
58363=>X"00",
58364=>X"00",
58365=>X"00",
58366=>X"00",
58367=>X"00",
58368=>X"00",
58369=>X"00",
58370=>X"00",
58371=>X"00",
58372=>X"00",
58373=>X"00",
58374=>X"00",
58375=>X"00",
58376=>X"00",
58377=>X"00",
58378=>X"00",
58379=>X"00",
58380=>X"00",
58381=>X"00",
58382=>X"00",
58383=>X"00",
58384=>X"00",
58385=>X"00",
58386=>X"00",
58387=>X"00",
58388=>X"00",
58389=>X"00",
58390=>X"00",
58391=>X"00",
58392=>X"00",
58393=>X"00",
58394=>X"00",
58395=>X"00",
58396=>X"00",
58397=>X"00",
58398=>X"00",
58399=>X"00",
58400=>X"00",
58401=>X"00",
58402=>X"00",
58403=>X"00",
58404=>X"00",
58405=>X"00",
58406=>X"00",
58407=>X"00",
58408=>X"00",
58409=>X"00",
58410=>X"00",
58411=>X"00",
58412=>X"00",
58413=>X"00",
58414=>X"00",
58415=>X"00",
58416=>X"00",
58417=>X"00",
58418=>X"00",
58419=>X"00",
58420=>X"00",
58421=>X"00",
58422=>X"00",
58423=>X"00",
58424=>X"00",
58425=>X"00",
58426=>X"00",
58427=>X"00",
58428=>X"00",
58429=>X"00",
58430=>X"00",
58431=>X"00",
58432=>X"00",
58433=>X"00",
58434=>X"00",
58435=>X"00",
58436=>X"00",
58437=>X"00",
58438=>X"00",
58439=>X"00",
58440=>X"00",
58441=>X"00",
58442=>X"00",
58443=>X"00",
58444=>X"00",
58445=>X"00",
58446=>X"00",
58447=>X"00",
58448=>X"00",
58449=>X"00",
58450=>X"00",
58451=>X"00",
58452=>X"00",
58453=>X"00",
58454=>X"00",
58455=>X"00",
58456=>X"00",
58457=>X"00",
58458=>X"00",
58459=>X"00",
58460=>X"00",
58461=>X"00",
58462=>X"00",
58463=>X"00",
58464=>X"00",
58465=>X"00",
58466=>X"00",
58467=>X"00",
58468=>X"00",
58469=>X"00",
58470=>X"00",
58471=>X"00",
58472=>X"00",
58473=>X"00",
58474=>X"00",
58475=>X"00",
58476=>X"00",
58477=>X"00",
58478=>X"00",
58479=>X"00",
58480=>X"00",
58481=>X"00",
58482=>X"00",
58483=>X"00",
58484=>X"00",
58485=>X"00",
58486=>X"00",
58487=>X"00",
58488=>X"00",
58489=>X"00",
58490=>X"00",
58491=>X"00",
58492=>X"00",
58493=>X"00",
58494=>X"00",
58495=>X"00",
58496=>X"00",
58497=>X"00",
58498=>X"00",
58499=>X"00",
58500=>X"00",
58501=>X"00",
58502=>X"00",
58503=>X"00",
58504=>X"00",
58505=>X"00",
58506=>X"00",
58507=>X"00",
58508=>X"00",
58509=>X"00",
58510=>X"00",
58511=>X"00",
58512=>X"00",
58513=>X"00",
58514=>X"00",
58515=>X"00",
58516=>X"00",
58517=>X"00",
58518=>X"00",
58519=>X"00",
58520=>X"00",
58521=>X"00",
58522=>X"00",
58523=>X"00",
58524=>X"00",
58525=>X"00",
58526=>X"00",
58527=>X"00",
58528=>X"00",
58529=>X"00",
58530=>X"00",
58531=>X"00",
58532=>X"00",
58533=>X"00",
58534=>X"00",
58535=>X"00",
58536=>X"00",
58537=>X"00",
58538=>X"00",
58539=>X"00",
58540=>X"00",
58541=>X"00",
58542=>X"00",
58543=>X"00",
58544=>X"00",
58545=>X"00",
58546=>X"00",
58547=>X"00",
58548=>X"00",
58549=>X"00",
58550=>X"00",
58551=>X"00",
58552=>X"00",
58553=>X"00",
58554=>X"00",
58555=>X"00",
58556=>X"00",
58557=>X"00",
58558=>X"00",
58559=>X"00",
58560=>X"00",
58561=>X"00",
58562=>X"00",
58563=>X"00",
58564=>X"00",
58565=>X"00",
58566=>X"00",
58567=>X"00",
58568=>X"00",
58569=>X"00",
58570=>X"00",
58571=>X"00",
58572=>X"00",
58573=>X"00",
58574=>X"00",
58575=>X"00",
58576=>X"00",
58577=>X"00",
58578=>X"00",
58579=>X"00",
58580=>X"00",
58581=>X"00",
58582=>X"00",
58583=>X"00",
58584=>X"00",
58585=>X"00",
58586=>X"00",
58587=>X"00",
58588=>X"00",
58589=>X"00",
58590=>X"00",
58591=>X"00",
58592=>X"00",
58593=>X"00",
58594=>X"00",
58595=>X"00",
58596=>X"00",
58597=>X"00",
58598=>X"00",
58599=>X"00",
58600=>X"00",
58601=>X"00",
58602=>X"00",
58603=>X"00",
58604=>X"00",
58605=>X"00",
58606=>X"00",
58607=>X"00",
58608=>X"00",
58609=>X"00",
58610=>X"00",
58611=>X"00",
58612=>X"00",
58613=>X"00",
58614=>X"00",
58615=>X"00",
58616=>X"00",
58617=>X"00",
58618=>X"00",
58619=>X"00",
58620=>X"00",
58621=>X"00",
58622=>X"00",
58623=>X"00",
58624=>X"00",
58625=>X"00",
58626=>X"00",
58627=>X"00",
58628=>X"00",
58629=>X"00",
58630=>X"00",
58631=>X"00",
58632=>X"00",
58633=>X"00",
58634=>X"00",
58635=>X"00",
58636=>X"00",
58637=>X"00",
58638=>X"00",
58639=>X"00",
58640=>X"00",
58641=>X"00",
58642=>X"00",
58643=>X"00",
58644=>X"00",
58645=>X"00",
58646=>X"00",
58647=>X"00",
58648=>X"00",
58649=>X"00",
58650=>X"00",
58651=>X"00",
58652=>X"00",
58653=>X"00",
58654=>X"00",
58655=>X"00",
58656=>X"00",
58657=>X"00",
58658=>X"00",
58659=>X"00",
58660=>X"00",
58661=>X"00",
58662=>X"00",
58663=>X"00",
58664=>X"00",
58665=>X"00",
58666=>X"00",
58667=>X"00",
58668=>X"00",
58669=>X"00",
58670=>X"00",
58671=>X"00",
58672=>X"00",
58673=>X"00",
58674=>X"00",
58675=>X"00",
58676=>X"00",
58677=>X"00",
58678=>X"00",
58679=>X"00",
58680=>X"00",
58681=>X"00",
58682=>X"00",
58683=>X"00",
58684=>X"00",
58685=>X"00",
58686=>X"00",
58687=>X"00",
58688=>X"00",
58689=>X"00",
58690=>X"00",
58691=>X"00",
58692=>X"00",
58693=>X"00",
58694=>X"00",
58695=>X"00",
58696=>X"00",
58697=>X"00",
58698=>X"00",
58699=>X"00",
58700=>X"00",
58701=>X"00",
58702=>X"00",
58703=>X"00",
58704=>X"00",
58705=>X"00",
58706=>X"00",
58707=>X"00",
58708=>X"00",
58709=>X"00",
58710=>X"00",
58711=>X"00",
58712=>X"00",
58713=>X"00",
58714=>X"00",
58715=>X"00",
58716=>X"00",
58717=>X"00",
58718=>X"00",
58719=>X"00",
58720=>X"00",
58721=>X"00",
58722=>X"00",
58723=>X"00",
58724=>X"00",
58725=>X"00",
58726=>X"00",
58727=>X"00",
58728=>X"00",
58729=>X"00",
58730=>X"00",
58731=>X"00",
58732=>X"00",
58733=>X"00",
58734=>X"00",
58735=>X"00",
58736=>X"00",
58737=>X"00",
58738=>X"00",
58739=>X"00",
58740=>X"00",
58741=>X"00",
58742=>X"00",
58743=>X"00",
58744=>X"00",
58745=>X"00",
58746=>X"00",
58747=>X"00",
58748=>X"00",
58749=>X"00",
58750=>X"00",
58751=>X"00",
58752=>X"00",
58753=>X"00",
58754=>X"00",
58755=>X"00",
58756=>X"00",
58757=>X"00",
58758=>X"00",
58759=>X"00",
58760=>X"00",
58761=>X"00",
58762=>X"00",
58763=>X"00",
58764=>X"00",
58765=>X"00",
58766=>X"00",
58767=>X"00",
58768=>X"00",
58769=>X"00",
58770=>X"00",
58771=>X"00",
58772=>X"00",
58773=>X"00",
58774=>X"00",
58775=>X"00",
58776=>X"00",
58777=>X"00",
58778=>X"00",
58779=>X"00",
58780=>X"00",
58781=>X"00",
58782=>X"00",
58783=>X"00",
58784=>X"00",
58785=>X"00",
58786=>X"00",
58787=>X"00",
58788=>X"00",
58789=>X"00",
58790=>X"00",
58791=>X"00",
58792=>X"00",
58793=>X"00",
58794=>X"00",
58795=>X"00",
58796=>X"00",
58797=>X"00",
58798=>X"00",
58799=>X"00",
58800=>X"00",
58801=>X"00",
58802=>X"00",
58803=>X"00",
58804=>X"00",
58805=>X"00",
58806=>X"00",
58807=>X"00",
58808=>X"00",
58809=>X"00",
58810=>X"00",
58811=>X"00",
58812=>X"00",
58813=>X"00",
58814=>X"00",
58815=>X"00",
58816=>X"00",
58817=>X"00",
58818=>X"00",
58819=>X"00",
58820=>X"00",
58821=>X"00",
58822=>X"00",
58823=>X"00",
58824=>X"00",
58825=>X"00",
58826=>X"00",
58827=>X"00",
58828=>X"00",
58829=>X"00",
58830=>X"00",
58831=>X"00",
58832=>X"00",
58833=>X"00",
58834=>X"00",
58835=>X"00",
58836=>X"00",
58837=>X"00",
58838=>X"00",
58839=>X"00",
58840=>X"00",
58841=>X"00",
58842=>X"00",
58843=>X"00",
58844=>X"00",
58845=>X"00",
58846=>X"00",
58847=>X"00",
58848=>X"00",
58849=>X"00",
58850=>X"00",
58851=>X"00",
58852=>X"00",
58853=>X"00",
58854=>X"00",
58855=>X"00",
58856=>X"00",
58857=>X"00",
58858=>X"00",
58859=>X"00",
58860=>X"00",
58861=>X"00",
58862=>X"00",
58863=>X"00",
58864=>X"00",
58865=>X"00",
58866=>X"00",
58867=>X"00",
58868=>X"00",
58869=>X"00",
58870=>X"00",
58871=>X"00",
58872=>X"00",
58873=>X"00",
58874=>X"00",
58875=>X"00",
58876=>X"00",
58877=>X"00",
58878=>X"00",
58879=>X"00",
58880=>X"00",
58881=>X"00",
58882=>X"00",
58883=>X"00",
58884=>X"00",
58885=>X"00",
58886=>X"00",
58887=>X"00",
58888=>X"00",
58889=>X"00",
58890=>X"00",
58891=>X"00",
58892=>X"00",
58893=>X"00",
58894=>X"00",
58895=>X"00",
58896=>X"00",
58897=>X"00",
58898=>X"00",
58899=>X"00",
58900=>X"00",
58901=>X"00",
58902=>X"00",
58903=>X"00",
58904=>X"00",
58905=>X"00",
58906=>X"00",
58907=>X"00",
58908=>X"00",
58909=>X"00",
58910=>X"00",
58911=>X"00",
58912=>X"00",
58913=>X"00",
58914=>X"00",
58915=>X"00",
58916=>X"00",
58917=>X"00",
58918=>X"00",
58919=>X"00",
58920=>X"00",
58921=>X"00",
58922=>X"00",
58923=>X"00",
58924=>X"00",
58925=>X"00",
58926=>X"00",
58927=>X"00",
58928=>X"00",
58929=>X"00",
58930=>X"00",
58931=>X"00",
58932=>X"00",
58933=>X"00",
58934=>X"00",
58935=>X"00",
58936=>X"00",
58937=>X"00",
58938=>X"00",
58939=>X"00",
58940=>X"00",
58941=>X"00",
58942=>X"00",
58943=>X"00",
58944=>X"00",
58945=>X"00",
58946=>X"00",
58947=>X"00",
58948=>X"00",
58949=>X"00",
58950=>X"00",
58951=>X"00",
58952=>X"00",
58953=>X"00",
58954=>X"00",
58955=>X"00",
58956=>X"00",
58957=>X"00",
58958=>X"00",
58959=>X"00",
58960=>X"00",
58961=>X"00",
58962=>X"00",
58963=>X"00",
58964=>X"00",
58965=>X"00",
58966=>X"00",
58967=>X"00",
58968=>X"00",
58969=>X"00",
58970=>X"00",
58971=>X"00",
58972=>X"00",
58973=>X"00",
58974=>X"00",
58975=>X"00",
58976=>X"00",
58977=>X"00",
58978=>X"00",
58979=>X"00",
58980=>X"00",
58981=>X"00",
58982=>X"00",
58983=>X"00",
58984=>X"00",
58985=>X"00",
58986=>X"00",
58987=>X"00",
58988=>X"00",
58989=>X"00",
58990=>X"00",
58991=>X"00",
58992=>X"00",
58993=>X"00",
58994=>X"00",
58995=>X"00",
58996=>X"00",
58997=>X"00",
58998=>X"00",
58999=>X"00",
59000=>X"00",
59001=>X"00",
59002=>X"00",
59003=>X"00",
59004=>X"00",
59005=>X"00",
59006=>X"00",
59007=>X"00",
59008=>X"00",
59009=>X"00",
59010=>X"00",
59011=>X"00",
59012=>X"00",
59013=>X"00",
59014=>X"00",
59015=>X"00",
59016=>X"00",
59017=>X"00",
59018=>X"00",
59019=>X"00",
59020=>X"00",
59021=>X"00",
59022=>X"00",
59023=>X"00",
59024=>X"00",
59025=>X"00",
59026=>X"00",
59027=>X"00",
59028=>X"00",
59029=>X"00",
59030=>X"00",
59031=>X"00",
59032=>X"00",
59033=>X"00",
59034=>X"00",
59035=>X"00",
59036=>X"00",
59037=>X"00",
59038=>X"00",
59039=>X"00",
59040=>X"00",
59041=>X"00",
59042=>X"00",
59043=>X"00",
59044=>X"00",
59045=>X"00",
59046=>X"00",
59047=>X"00",
59048=>X"00",
59049=>X"00",
59050=>X"00",
59051=>X"00",
59052=>X"00",
59053=>X"00",
59054=>X"00",
59055=>X"00",
59056=>X"00",
59057=>X"00",
59058=>X"00",
59059=>X"00",
59060=>X"00",
59061=>X"00",
59062=>X"00",
59063=>X"00",
59064=>X"00",
59065=>X"00",
59066=>X"00",
59067=>X"00",
59068=>X"00",
59069=>X"00",
59070=>X"00",
59071=>X"00",
59072=>X"00",
59073=>X"00",
59074=>X"00",
59075=>X"00",
59076=>X"00",
59077=>X"00",
59078=>X"00",
59079=>X"00",
59080=>X"00",
59081=>X"00",
59082=>X"00",
59083=>X"00",
59084=>X"00",
59085=>X"00",
59086=>X"00",
59087=>X"00",
59088=>X"00",
59089=>X"00",
59090=>X"00",
59091=>X"00",
59092=>X"00",
59093=>X"00",
59094=>X"00",
59095=>X"00",
59096=>X"00",
59097=>X"00",
59098=>X"00",
59099=>X"00",
59100=>X"00",
59101=>X"00",
59102=>X"00",
59103=>X"00",
59104=>X"00",
59105=>X"00",
59106=>X"00",
59107=>X"00",
59108=>X"00",
59109=>X"00",
59110=>X"00",
59111=>X"00",
59112=>X"00",
59113=>X"00",
59114=>X"00",
59115=>X"00",
59116=>X"00",
59117=>X"00",
59118=>X"00",
59119=>X"00",
59120=>X"00",
59121=>X"00",
59122=>X"00",
59123=>X"00",
59124=>X"00",
59125=>X"00",
59126=>X"00",
59127=>X"00",
59128=>X"00",
59129=>X"00",
59130=>X"00",
59131=>X"00",
59132=>X"00",
59133=>X"00",
59134=>X"00",
59135=>X"00",
59136=>X"00",
59137=>X"00",
59138=>X"00",
59139=>X"00",
59140=>X"00",
59141=>X"00",
59142=>X"00",
59143=>X"00",
59144=>X"00",
59145=>X"00",
59146=>X"00",
59147=>X"00",
59148=>X"00",
59149=>X"00",
59150=>X"00",
59151=>X"00",
59152=>X"00",
59153=>X"00",
59154=>X"00",
59155=>X"00",
59156=>X"00",
59157=>X"00",
59158=>X"00",
59159=>X"00",
59160=>X"00",
59161=>X"00",
59162=>X"00",
59163=>X"00",
59164=>X"00",
59165=>X"00",
59166=>X"00",
59167=>X"00",
59168=>X"00",
59169=>X"00",
59170=>X"00",
59171=>X"00",
59172=>X"00",
59173=>X"00",
59174=>X"00",
59175=>X"00",
59176=>X"00",
59177=>X"00",
59178=>X"00",
59179=>X"00",
59180=>X"00",
59181=>X"00",
59182=>X"00",
59183=>X"00",
59184=>X"00",
59185=>X"00",
59186=>X"00",
59187=>X"00",
59188=>X"00",
59189=>X"00",
59190=>X"00",
59191=>X"00",
59192=>X"00",
59193=>X"00",
59194=>X"00",
59195=>X"00",
59196=>X"00",
59197=>X"00",
59198=>X"00",
59199=>X"00",
59200=>X"00",
59201=>X"00",
59202=>X"00",
59203=>X"00",
59204=>X"00",
59205=>X"00",
59206=>X"00",
59207=>X"00",
59208=>X"00",
59209=>X"00",
59210=>X"00",
59211=>X"00",
59212=>X"00",
59213=>X"00",
59214=>X"00",
59215=>X"00",
59216=>X"00",
59217=>X"00",
59218=>X"00",
59219=>X"00",
59220=>X"00",
59221=>X"00",
59222=>X"00",
59223=>X"00",
59224=>X"00",
59225=>X"00",
59226=>X"00",
59227=>X"00",
59228=>X"00",
59229=>X"00",
59230=>X"00",
59231=>X"00",
59232=>X"00",
59233=>X"00",
59234=>X"00",
59235=>X"00",
59236=>X"00",
59237=>X"00",
59238=>X"00",
59239=>X"00",
59240=>X"00",
59241=>X"00",
59242=>X"00",
59243=>X"00",
59244=>X"00",
59245=>X"00",
59246=>X"00",
59247=>X"00",
59248=>X"00",
59249=>X"00",
59250=>X"00",
59251=>X"00",
59252=>X"00",
59253=>X"00",
59254=>X"00",
59255=>X"00",
59256=>X"00",
59257=>X"00",
59258=>X"00",
59259=>X"00",
59260=>X"00",
59261=>X"00",
59262=>X"00",
59263=>X"00",
59264=>X"00",
59265=>X"00",
59266=>X"00",
59267=>X"00",
59268=>X"00",
59269=>X"00",
59270=>X"00",
59271=>X"00",
59272=>X"00",
59273=>X"00",
59274=>X"00",
59275=>X"00",
59276=>X"00",
59277=>X"00",
59278=>X"00",
59279=>X"00",
59280=>X"00",
59281=>X"00",
59282=>X"00",
59283=>X"00",
59284=>X"00",
59285=>X"00",
59286=>X"00",
59287=>X"00",
59288=>X"00",
59289=>X"00",
59290=>X"00",
59291=>X"00",
59292=>X"00",
59293=>X"00",
59294=>X"00",
59295=>X"00",
59296=>X"00",
59297=>X"00",
59298=>X"00",
59299=>X"00",
59300=>X"00",
59301=>X"00",
59302=>X"00",
59303=>X"00",
59304=>X"00",
59305=>X"00",
59306=>X"00",
59307=>X"00",
59308=>X"00",
59309=>X"00",
59310=>X"00",
59311=>X"00",
59312=>X"00",
59313=>X"00",
59314=>X"00",
59315=>X"00",
59316=>X"00",
59317=>X"00",
59318=>X"00",
59319=>X"00",
59320=>X"00",
59321=>X"00",
59322=>X"00",
59323=>X"00",
59324=>X"00",
59325=>X"00",
59326=>X"00",
59327=>X"00",
59328=>X"00",
59329=>X"00",
59330=>X"00",
59331=>X"00",
59332=>X"00",
59333=>X"00",
59334=>X"00",
59335=>X"00",
59336=>X"00",
59337=>X"00",
59338=>X"00",
59339=>X"00",
59340=>X"00",
59341=>X"00",
59342=>X"00",
59343=>X"00",
59344=>X"00",
59345=>X"00",
59346=>X"00",
59347=>X"00",
59348=>X"00",
59349=>X"00",
59350=>X"00",
59351=>X"00",
59352=>X"00",
59353=>X"00",
59354=>X"00",
59355=>X"00",
59356=>X"00",
59357=>X"00",
59358=>X"00",
59359=>X"00",
59360=>X"00",
59361=>X"00",
59362=>X"00",
59363=>X"00",
59364=>X"00",
59365=>X"00",
59366=>X"00",
59367=>X"00",
59368=>X"00",
59369=>X"00",
59370=>X"00",
59371=>X"00",
59372=>X"00",
59373=>X"00",
59374=>X"00",
59375=>X"00",
59376=>X"00",
59377=>X"00",
59378=>X"00",
59379=>X"00",
59380=>X"00",
59381=>X"00",
59382=>X"00",
59383=>X"00",
59384=>X"00",
59385=>X"00",
59386=>X"00",
59387=>X"00",
59388=>X"00",
59389=>X"00",
59390=>X"00",
59391=>X"00",
59392=>X"00",
59393=>X"00",
59394=>X"00",
59395=>X"00",
59396=>X"00",
59397=>X"00",
59398=>X"00",
59399=>X"00",
59400=>X"00",
59401=>X"00",
59402=>X"00",
59403=>X"00",
59404=>X"00",
59405=>X"00",
59406=>X"00",
59407=>X"00",
59408=>X"00",
59409=>X"00",
59410=>X"00",
59411=>X"00",
59412=>X"00",
59413=>X"00",
59414=>X"00",
59415=>X"00",
59416=>X"00",
59417=>X"00",
59418=>X"00",
59419=>X"00",
59420=>X"00",
59421=>X"00",
59422=>X"00",
59423=>X"00",
59424=>X"00",
59425=>X"00",
59426=>X"00",
59427=>X"00",
59428=>X"00",
59429=>X"00",
59430=>X"00",
59431=>X"00",
59432=>X"00",
59433=>X"00",
59434=>X"00",
59435=>X"00",
59436=>X"00",
59437=>X"00",
59438=>X"00",
59439=>X"00",
59440=>X"00",
59441=>X"00",
59442=>X"00",
59443=>X"00",
59444=>X"00",
59445=>X"00",
59446=>X"00",
59447=>X"00",
59448=>X"00",
59449=>X"00",
59450=>X"00",
59451=>X"00",
59452=>X"00",
59453=>X"00",
59454=>X"00",
59455=>X"00",
59456=>X"00",
59457=>X"00",
59458=>X"00",
59459=>X"00",
59460=>X"00",
59461=>X"00",
59462=>X"00",
59463=>X"00",
59464=>X"00",
59465=>X"00",
59466=>X"00",
59467=>X"00",
59468=>X"00",
59469=>X"00",
59470=>X"00",
59471=>X"00",
59472=>X"00",
59473=>X"00",
59474=>X"00",
59475=>X"00",
59476=>X"00",
59477=>X"00",
59478=>X"00",
59479=>X"00",
59480=>X"00",
59481=>X"00",
59482=>X"00",
59483=>X"00",
59484=>X"00",
59485=>X"00",
59486=>X"00",
59487=>X"00",
59488=>X"00",
59489=>X"00",
59490=>X"00",
59491=>X"00",
59492=>X"00",
59493=>X"00",
59494=>X"00",
59495=>X"00",
59496=>X"00",
59497=>X"00",
59498=>X"00",
59499=>X"00",
59500=>X"00",
59501=>X"00",
59502=>X"00",
59503=>X"00",
59504=>X"00",
59505=>X"00",
59506=>X"00",
59507=>X"00",
59508=>X"00",
59509=>X"00",
59510=>X"00",
59511=>X"00",
59512=>X"00",
59513=>X"00",
59514=>X"00",
59515=>X"00",
59516=>X"00",
59517=>X"00",
59518=>X"00",
59519=>X"00",
59520=>X"00",
59521=>X"00",
59522=>X"00",
59523=>X"00",
59524=>X"00",
59525=>X"00",
59526=>X"00",
59527=>X"00",
59528=>X"00",
59529=>X"00",
59530=>X"00",
59531=>X"00",
59532=>X"00",
59533=>X"00",
59534=>X"00",
59535=>X"00",
59536=>X"00",
59537=>X"00",
59538=>X"00",
59539=>X"00",
59540=>X"00",
59541=>X"00",
59542=>X"00",
59543=>X"00",
59544=>X"00",
59545=>X"00",
59546=>X"00",
59547=>X"00",
59548=>X"00",
59549=>X"00",
59550=>X"00",
59551=>X"00",
59552=>X"00",
59553=>X"00",
59554=>X"00",
59555=>X"00",
59556=>X"00",
59557=>X"00",
59558=>X"00",
59559=>X"00",
59560=>X"00",
59561=>X"00",
59562=>X"00",
59563=>X"00",
59564=>X"00",
59565=>X"00",
59566=>X"00",
59567=>X"00",
59568=>X"00",
59569=>X"00",
59570=>X"00",
59571=>X"00",
59572=>X"00",
59573=>X"00",
59574=>X"00",
59575=>X"00",
59576=>X"00",
59577=>X"00",
59578=>X"00",
59579=>X"00",
59580=>X"00",
59581=>X"00",
59582=>X"00",
59583=>X"00",
59584=>X"00",
59585=>X"00",
59586=>X"00",
59587=>X"00",
59588=>X"00",
59589=>X"00",
59590=>X"00",
59591=>X"00",
59592=>X"00",
59593=>X"00",
59594=>X"00",
59595=>X"00",
59596=>X"00",
59597=>X"00",
59598=>X"00",
59599=>X"00",
59600=>X"00",
59601=>X"00",
59602=>X"00",
59603=>X"00",
59604=>X"00",
59605=>X"00",
59606=>X"00",
59607=>X"00",
59608=>X"00",
59609=>X"00",
59610=>X"00",
59611=>X"00",
59612=>X"00",
59613=>X"00",
59614=>X"00",
59615=>X"00",
59616=>X"00",
59617=>X"00",
59618=>X"00",
59619=>X"00",
59620=>X"00",
59621=>X"00",
59622=>X"00",
59623=>X"00",
59624=>X"00",
59625=>X"00",
59626=>X"00",
59627=>X"00",
59628=>X"00",
59629=>X"00",
59630=>X"00",
59631=>X"00",
59632=>X"00",
59633=>X"00",
59634=>X"00",
59635=>X"00",
59636=>X"00",
59637=>X"00",
59638=>X"00",
59639=>X"00",
59640=>X"00",
59641=>X"00",
59642=>X"00",
59643=>X"00",
59644=>X"00",
59645=>X"00",
59646=>X"00",
59647=>X"00",
59648=>X"00",
59649=>X"00",
59650=>X"00",
59651=>X"00",
59652=>X"00",
59653=>X"00",
59654=>X"00",
59655=>X"00",
59656=>X"00",
59657=>X"00",
59658=>X"00",
59659=>X"00",
59660=>X"00",
59661=>X"00",
59662=>X"00",
59663=>X"00",
59664=>X"00",
59665=>X"00",
59666=>X"00",
59667=>X"00",
59668=>X"00",
59669=>X"00",
59670=>X"00",
59671=>X"00",
59672=>X"00",
59673=>X"00",
59674=>X"00",
59675=>X"00",
59676=>X"00",
59677=>X"00",
59678=>X"00",
59679=>X"00",
59680=>X"00",
59681=>X"00",
59682=>X"00",
59683=>X"00",
59684=>X"00",
59685=>X"00",
59686=>X"00",
59687=>X"00",
59688=>X"00",
59689=>X"00",
59690=>X"00",
59691=>X"00",
59692=>X"00",
59693=>X"00",
59694=>X"00",
59695=>X"00",
59696=>X"00",
59697=>X"00",
59698=>X"00",
59699=>X"00",
59700=>X"00",
59701=>X"00",
59702=>X"00",
59703=>X"00",
59704=>X"00",
59705=>X"00",
59706=>X"00",
59707=>X"00",
59708=>X"00",
59709=>X"00",
59710=>X"00",
59711=>X"00",
59712=>X"00",
59713=>X"00",
59714=>X"00",
59715=>X"00",
59716=>X"00",
59717=>X"00",
59718=>X"00",
59719=>X"00",
59720=>X"00",
59721=>X"00",
59722=>X"00",
59723=>X"00",
59724=>X"00",
59725=>X"00",
59726=>X"00",
59727=>X"00",
59728=>X"00",
59729=>X"00",
59730=>X"00",
59731=>X"00",
59732=>X"00",
59733=>X"00",
59734=>X"00",
59735=>X"00",
59736=>X"00",
59737=>X"00",
59738=>X"00",
59739=>X"00",
59740=>X"00",
59741=>X"00",
59742=>X"00",
59743=>X"00",
59744=>X"00",
59745=>X"00",
59746=>X"00",
59747=>X"00",
59748=>X"00",
59749=>X"00",
59750=>X"00",
59751=>X"00",
59752=>X"00",
59753=>X"00",
59754=>X"00",
59755=>X"00",
59756=>X"00",
59757=>X"00",
59758=>X"00",
59759=>X"00",
59760=>X"00",
59761=>X"00",
59762=>X"00",
59763=>X"00",
59764=>X"00",
59765=>X"00",
59766=>X"00",
59767=>X"00",
59768=>X"00",
59769=>X"00",
59770=>X"00",
59771=>X"00",
59772=>X"00",
59773=>X"00",
59774=>X"00",
59775=>X"00",
59776=>X"00",
59777=>X"00",
59778=>X"00",
59779=>X"00",
59780=>X"00",
59781=>X"00",
59782=>X"00",
59783=>X"00",
59784=>X"00",
59785=>X"00",
59786=>X"00",
59787=>X"00",
59788=>X"00",
59789=>X"00",
59790=>X"00",
59791=>X"00",
59792=>X"00",
59793=>X"00",
59794=>X"00",
59795=>X"00",
59796=>X"00",
59797=>X"00",
59798=>X"00",
59799=>X"00",
59800=>X"00",
59801=>X"00",
59802=>X"00",
59803=>X"00",
59804=>X"00",
59805=>X"00",
59806=>X"00",
59807=>X"00",
59808=>X"00",
59809=>X"00",
59810=>X"00",
59811=>X"00",
59812=>X"00",
59813=>X"00",
59814=>X"00",
59815=>X"00",
59816=>X"00",
59817=>X"00",
59818=>X"00",
59819=>X"00",
59820=>X"00",
59821=>X"00",
59822=>X"00",
59823=>X"00",
59824=>X"00",
59825=>X"00",
59826=>X"00",
59827=>X"00",
59828=>X"00",
59829=>X"00",
59830=>X"00",
59831=>X"00",
59832=>X"00",
59833=>X"00",
59834=>X"00",
59835=>X"00",
59836=>X"00",
59837=>X"00",
59838=>X"00",
59839=>X"00",
59840=>X"00",
59841=>X"00",
59842=>X"00",
59843=>X"00",
59844=>X"00",
59845=>X"00",
59846=>X"00",
59847=>X"00",
59848=>X"00",
59849=>X"00",
59850=>X"00",
59851=>X"00",
59852=>X"00",
59853=>X"00",
59854=>X"00",
59855=>X"00",
59856=>X"00",
59857=>X"00",
59858=>X"00",
59859=>X"00",
59860=>X"00",
59861=>X"00",
59862=>X"00",
59863=>X"00",
59864=>X"00",
59865=>X"00",
59866=>X"00",
59867=>X"00",
59868=>X"00",
59869=>X"00",
59870=>X"00",
59871=>X"00",
59872=>X"00",
59873=>X"00",
59874=>X"00",
59875=>X"00",
59876=>X"00",
59877=>X"00",
59878=>X"00",
59879=>X"00",
59880=>X"00",
59881=>X"00",
59882=>X"00",
59883=>X"00",
59884=>X"00",
59885=>X"00",
59886=>X"00",
59887=>X"00",
59888=>X"00",
59889=>X"00",
59890=>X"00",
59891=>X"00",
59892=>X"00",
59893=>X"00",
59894=>X"00",
59895=>X"00",
59896=>X"00",
59897=>X"00",
59898=>X"00",
59899=>X"00",
59900=>X"00",
59901=>X"00",
59902=>X"00",
59903=>X"00",
59904=>X"00",
59905=>X"00",
59906=>X"00",
59907=>X"00",
59908=>X"00",
59909=>X"00",
59910=>X"00",
59911=>X"00",
59912=>X"00",
59913=>X"00",
59914=>X"00",
59915=>X"00",
59916=>X"00",
59917=>X"00",
59918=>X"00",
59919=>X"00",
59920=>X"00",
59921=>X"00",
59922=>X"00",
59923=>X"00",
59924=>X"00",
59925=>X"00",
59926=>X"00",
59927=>X"00",
59928=>X"00",
59929=>X"00",
59930=>X"00",
59931=>X"00",
59932=>X"00",
59933=>X"00",
59934=>X"00",
59935=>X"00",
59936=>X"00",
59937=>X"00",
59938=>X"00",
59939=>X"00",
59940=>X"00",
59941=>X"00",
59942=>X"00",
59943=>X"00",
59944=>X"00",
59945=>X"00",
59946=>X"00",
59947=>X"00",
59948=>X"00",
59949=>X"00",
59950=>X"00",
59951=>X"00",
59952=>X"00",
59953=>X"00",
59954=>X"00",
59955=>X"00",
59956=>X"00",
59957=>X"00",
59958=>X"00",
59959=>X"00",
59960=>X"00",
59961=>X"00",
59962=>X"00",
59963=>X"00",
59964=>X"00",
59965=>X"00",
59966=>X"00",
59967=>X"00",
59968=>X"00",
59969=>X"00",
59970=>X"00",
59971=>X"00",
59972=>X"00",
59973=>X"00",
59974=>X"00",
59975=>X"00",
59976=>X"00",
59977=>X"00",
59978=>X"00",
59979=>X"00",
59980=>X"00",
59981=>X"00",
59982=>X"00",
59983=>X"00",
59984=>X"00",
59985=>X"00",
59986=>X"00",
59987=>X"00",
59988=>X"00",
59989=>X"00",
59990=>X"00",
59991=>X"00",
59992=>X"00",
59993=>X"00",
59994=>X"00",
59995=>X"00",
59996=>X"00",
59997=>X"00",
59998=>X"00",
59999=>X"00",
60000=>X"00",
60001=>X"00",
60002=>X"00",
60003=>X"00",
60004=>X"00",
60005=>X"00",
60006=>X"00",
60007=>X"00",
60008=>X"00",
60009=>X"00",
60010=>X"00",
60011=>X"00",
60012=>X"00",
60013=>X"00",
60014=>X"00",
60015=>X"00",
60016=>X"00",
60017=>X"00",
60018=>X"00",
60019=>X"00",
60020=>X"00",
60021=>X"00",
60022=>X"00",
60023=>X"00",
60024=>X"00",
60025=>X"00",
60026=>X"00",
60027=>X"00",
60028=>X"00",
60029=>X"00",
60030=>X"00",
60031=>X"00",
60032=>X"00",
60033=>X"00",
60034=>X"00",
60035=>X"00",
60036=>X"00",
60037=>X"00",
60038=>X"00",
60039=>X"00",
60040=>X"00",
60041=>X"00",
60042=>X"00",
60043=>X"00",
60044=>X"00",
60045=>X"00",
60046=>X"00",
60047=>X"00",
60048=>X"00",
60049=>X"00",
60050=>X"00",
60051=>X"00",
60052=>X"00",
60053=>X"00",
60054=>X"00",
60055=>X"00",
60056=>X"00",
60057=>X"00",
60058=>X"00",
60059=>X"00",
60060=>X"00",
60061=>X"00",
60062=>X"00",
60063=>X"00",
60064=>X"00",
60065=>X"00",
60066=>X"00",
60067=>X"00",
60068=>X"00",
60069=>X"00",
60070=>X"00",
60071=>X"00",
60072=>X"00",
60073=>X"00",
60074=>X"00",
60075=>X"00",
60076=>X"00",
60077=>X"00",
60078=>X"00",
60079=>X"00",
60080=>X"00",
60081=>X"00",
60082=>X"00",
60083=>X"00",
60084=>X"00",
60085=>X"00",
60086=>X"00",
60087=>X"00",
60088=>X"00",
60089=>X"00",
60090=>X"00",
60091=>X"00",
60092=>X"00",
60093=>X"00",
60094=>X"00",
60095=>X"00",
60096=>X"00",
60097=>X"00",
60098=>X"00",
60099=>X"00",
60100=>X"00",
60101=>X"00",
60102=>X"00",
60103=>X"00",
60104=>X"00",
60105=>X"00",
60106=>X"00",
60107=>X"00",
60108=>X"00",
60109=>X"00",
60110=>X"00",
60111=>X"00",
60112=>X"00",
60113=>X"00",
60114=>X"00",
60115=>X"00",
60116=>X"00",
60117=>X"00",
60118=>X"00",
60119=>X"00",
60120=>X"00",
60121=>X"00",
60122=>X"00",
60123=>X"00",
60124=>X"00",
60125=>X"00",
60126=>X"00",
60127=>X"00",
60128=>X"00",
60129=>X"00",
60130=>X"00",
60131=>X"00",
60132=>X"00",
60133=>X"00",
60134=>X"00",
60135=>X"00",
60136=>X"00",
60137=>X"00",
60138=>X"00",
60139=>X"00",
60140=>X"00",
60141=>X"00",
60142=>X"00",
60143=>X"00",
60144=>X"00",
60145=>X"00",
60146=>X"00",
60147=>X"00",
60148=>X"00",
60149=>X"00",
60150=>X"00",
60151=>X"00",
60152=>X"00",
60153=>X"00",
60154=>X"00",
60155=>X"00",
60156=>X"00",
60157=>X"00",
60158=>X"00",
60159=>X"00",
60160=>X"00",
60161=>X"00",
60162=>X"00",
60163=>X"00",
60164=>X"00",
60165=>X"00",
60166=>X"00",
60167=>X"00",
60168=>X"00",
60169=>X"00",
60170=>X"00",
60171=>X"00",
60172=>X"00",
60173=>X"00",
60174=>X"00",
60175=>X"00",
60176=>X"00",
60177=>X"00",
60178=>X"00",
60179=>X"00",
60180=>X"00",
60181=>X"00",
60182=>X"00",
60183=>X"00",
60184=>X"00",
60185=>X"00",
60186=>X"00",
60187=>X"00",
60188=>X"00",
60189=>X"00",
60190=>X"00",
60191=>X"00",
60192=>X"00",
60193=>X"00",
60194=>X"00",
60195=>X"00",
60196=>X"00",
60197=>X"00",
60198=>X"00",
60199=>X"00",
60200=>X"00",
60201=>X"00",
60202=>X"00",
60203=>X"00",
60204=>X"00",
60205=>X"00",
60206=>X"00",
60207=>X"00",
60208=>X"00",
60209=>X"00",
60210=>X"00",
60211=>X"00",
60212=>X"00",
60213=>X"00",
60214=>X"00",
60215=>X"00",
60216=>X"00",
60217=>X"00",
60218=>X"00",
60219=>X"00",
60220=>X"00",
60221=>X"00",
60222=>X"00",
60223=>X"00",
60224=>X"00",
60225=>X"00",
60226=>X"00",
60227=>X"00",
60228=>X"00",
60229=>X"00",
60230=>X"00",
60231=>X"00",
60232=>X"00",
60233=>X"00",
60234=>X"00",
60235=>X"00",
60236=>X"00",
60237=>X"00",
60238=>X"00",
60239=>X"00",
60240=>X"00",
60241=>X"00",
60242=>X"00",
60243=>X"00",
60244=>X"00",
60245=>X"00",
60246=>X"00",
60247=>X"00",
60248=>X"00",
60249=>X"00",
60250=>X"00",
60251=>X"00",
60252=>X"00",
60253=>X"00",
60254=>X"00",
60255=>X"00",
60256=>X"00",
60257=>X"00",
60258=>X"00",
60259=>X"00",
60260=>X"00",
60261=>X"00",
60262=>X"00",
60263=>X"00",
60264=>X"00",
60265=>X"00",
60266=>X"00",
60267=>X"00",
60268=>X"00",
60269=>X"00",
60270=>X"00",
60271=>X"00",
60272=>X"00",
60273=>X"00",
60274=>X"00",
60275=>X"00",
60276=>X"00",
60277=>X"00",
60278=>X"00",
60279=>X"00",
60280=>X"00",
60281=>X"00",
60282=>X"00",
60283=>X"00",
60284=>X"00",
60285=>X"00",
60286=>X"00",
60287=>X"00",
60288=>X"00",
60289=>X"00",
60290=>X"00",
60291=>X"00",
60292=>X"00",
60293=>X"00",
60294=>X"00",
60295=>X"00",
60296=>X"00",
60297=>X"00",
60298=>X"00",
60299=>X"00",
60300=>X"00",
60301=>X"00",
60302=>X"00",
60303=>X"00",
60304=>X"00",
60305=>X"00",
60306=>X"00",
60307=>X"00",
60308=>X"00",
60309=>X"00",
60310=>X"00",
60311=>X"00",
60312=>X"00",
60313=>X"00",
60314=>X"00",
60315=>X"00",
60316=>X"00",
60317=>X"00",
60318=>X"00",
60319=>X"00",
60320=>X"00",
60321=>X"00",
60322=>X"00",
60323=>X"00",
60324=>X"00",
60325=>X"00",
60326=>X"00",
60327=>X"00",
60328=>X"00",
60329=>X"00",
60330=>X"00",
60331=>X"00",
60332=>X"00",
60333=>X"00",
60334=>X"00",
60335=>X"00",
60336=>X"00",
60337=>X"00",
60338=>X"00",
60339=>X"00",
60340=>X"00",
60341=>X"00",
60342=>X"00",
60343=>X"00",
60344=>X"00",
60345=>X"00",
60346=>X"00",
60347=>X"00",
60348=>X"00",
60349=>X"00",
60350=>X"00",
60351=>X"00",
60352=>X"00",
60353=>X"00",
60354=>X"00",
60355=>X"00",
60356=>X"00",
60357=>X"00",
60358=>X"00",
60359=>X"00",
60360=>X"00",
60361=>X"00",
60362=>X"00",
60363=>X"00",
60364=>X"00",
60365=>X"00",
60366=>X"00",
60367=>X"00",
60368=>X"00",
60369=>X"00",
60370=>X"00",
60371=>X"00",
60372=>X"00",
60373=>X"00",
60374=>X"00",
60375=>X"00",
60376=>X"00",
60377=>X"00",
60378=>X"00",
60379=>X"00",
60380=>X"00",
60381=>X"00",
60382=>X"00",
60383=>X"00",
60384=>X"00",
60385=>X"00",
60386=>X"00",
60387=>X"00",
60388=>X"00",
60389=>X"00",
60390=>X"00",
60391=>X"00",
60392=>X"00",
60393=>X"00",
60394=>X"00",
60395=>X"00",
60396=>X"00",
60397=>X"00",
60398=>X"00",
60399=>X"00",
60400=>X"00",
60401=>X"00",
60402=>X"00",
60403=>X"00",
60404=>X"00",
60405=>X"00",
60406=>X"00",
60407=>X"00",
60408=>X"00",
60409=>X"00",
60410=>X"00",
60411=>X"00",
60412=>X"00",
60413=>X"00",
60414=>X"00",
60415=>X"00",
60416=>X"00",
60417=>X"00",
60418=>X"00",
60419=>X"00",
60420=>X"00",
60421=>X"00",
60422=>X"00",
60423=>X"00",
60424=>X"00",
60425=>X"00",
60426=>X"00",
60427=>X"00",
60428=>X"00",
60429=>X"00",
60430=>X"00",
60431=>X"00",
60432=>X"00",
60433=>X"00",
60434=>X"00",
60435=>X"00",
60436=>X"00",
60437=>X"00",
60438=>X"00",
60439=>X"00",
60440=>X"00",
60441=>X"00",
60442=>X"00",
60443=>X"00",
60444=>X"00",
60445=>X"00",
60446=>X"00",
60447=>X"00",
60448=>X"00",
60449=>X"00",
60450=>X"00",
60451=>X"00",
60452=>X"00",
60453=>X"00",
60454=>X"00",
60455=>X"00",
60456=>X"00",
60457=>X"00",
60458=>X"00",
60459=>X"00",
60460=>X"00",
60461=>X"00",
60462=>X"00",
60463=>X"00",
60464=>X"00",
60465=>X"00",
60466=>X"00",
60467=>X"00",
60468=>X"00",
60469=>X"00",
60470=>X"00",
60471=>X"00",
60472=>X"00",
60473=>X"00",
60474=>X"00",
60475=>X"00",
60476=>X"00",
60477=>X"00",
60478=>X"00",
60479=>X"00",
60480=>X"00",
60481=>X"00",
60482=>X"00",
60483=>X"00",
60484=>X"00",
60485=>X"00",
60486=>X"00",
60487=>X"00",
60488=>X"00",
60489=>X"00",
60490=>X"00",
60491=>X"00",
60492=>X"00",
60493=>X"00",
60494=>X"00",
60495=>X"00",
60496=>X"00",
60497=>X"00",
60498=>X"00",
60499=>X"00",
60500=>X"00",
60501=>X"00",
60502=>X"00",
60503=>X"00",
60504=>X"00",
60505=>X"00",
60506=>X"00",
60507=>X"00",
60508=>X"00",
60509=>X"00",
60510=>X"00",
60511=>X"00",
60512=>X"00",
60513=>X"00",
60514=>X"00",
60515=>X"00",
60516=>X"00",
60517=>X"00",
60518=>X"00",
60519=>X"00",
60520=>X"00",
60521=>X"00",
60522=>X"00",
60523=>X"00",
60524=>X"00",
60525=>X"00",
60526=>X"00",
60527=>X"00",
60528=>X"00",
60529=>X"00",
60530=>X"00",
60531=>X"00",
60532=>X"00",
60533=>X"00",
60534=>X"00",
60535=>X"00",
60536=>X"00",
60537=>X"00",
60538=>X"00",
60539=>X"00",
60540=>X"00",
60541=>X"00",
60542=>X"00",
60543=>X"00",
60544=>X"00",
60545=>X"00",
60546=>X"00",
60547=>X"00",
60548=>X"00",
60549=>X"00",
60550=>X"00",
60551=>X"00",
60552=>X"00",
60553=>X"00",
60554=>X"00",
60555=>X"00",
60556=>X"00",
60557=>X"00",
60558=>X"00",
60559=>X"00",
60560=>X"00",
60561=>X"00",
60562=>X"00",
60563=>X"00",
60564=>X"00",
60565=>X"00",
60566=>X"00",
60567=>X"00",
60568=>X"00",
60569=>X"00",
60570=>X"00",
60571=>X"00",
60572=>X"00",
60573=>X"00",
60574=>X"00",
60575=>X"00",
60576=>X"00",
60577=>X"00",
60578=>X"00",
60579=>X"00",
60580=>X"00",
60581=>X"00",
60582=>X"00",
60583=>X"00",
60584=>X"00",
60585=>X"00",
60586=>X"00",
60587=>X"00",
60588=>X"00",
60589=>X"00",
60590=>X"00",
60591=>X"00",
60592=>X"00",
60593=>X"00",
60594=>X"00",
60595=>X"00",
60596=>X"00",
60597=>X"00",
60598=>X"00",
60599=>X"00",
60600=>X"00",
60601=>X"00",
60602=>X"00",
60603=>X"00",
60604=>X"00",
60605=>X"00",
60606=>X"00",
60607=>X"00",
60608=>X"00",
60609=>X"00",
60610=>X"00",
60611=>X"00",
60612=>X"00",
60613=>X"00",
60614=>X"00",
60615=>X"00",
60616=>X"00",
60617=>X"00",
60618=>X"00",
60619=>X"00",
60620=>X"00",
60621=>X"00",
60622=>X"00",
60623=>X"00",
60624=>X"00",
60625=>X"00",
60626=>X"00",
60627=>X"00",
60628=>X"00",
60629=>X"00",
60630=>X"00",
60631=>X"00",
60632=>X"00",
60633=>X"00",
60634=>X"00",
60635=>X"00",
60636=>X"00",
60637=>X"00",
60638=>X"00",
60639=>X"00",
60640=>X"00",
60641=>X"00",
60642=>X"00",
60643=>X"00",
60644=>X"00",
60645=>X"00",
60646=>X"00",
60647=>X"00",
60648=>X"00",
60649=>X"00",
60650=>X"00",
60651=>X"00",
60652=>X"00",
60653=>X"00",
60654=>X"00",
60655=>X"00",
60656=>X"00",
60657=>X"00",
60658=>X"00",
60659=>X"00",
60660=>X"00",
60661=>X"00",
60662=>X"00",
60663=>X"00",
60664=>X"00",
60665=>X"00",
60666=>X"00",
60667=>X"00",
60668=>X"00",
60669=>X"00",
60670=>X"00",
60671=>X"00",
60672=>X"00",
60673=>X"00",
60674=>X"00",
60675=>X"00",
60676=>X"00",
60677=>X"00",
60678=>X"00",
60679=>X"00",
60680=>X"00",
60681=>X"00",
60682=>X"00",
60683=>X"00",
60684=>X"00",
60685=>X"00",
60686=>X"00",
60687=>X"00",
60688=>X"00",
60689=>X"00",
60690=>X"00",
60691=>X"00",
60692=>X"00",
60693=>X"00",
60694=>X"00",
60695=>X"00",
60696=>X"00",
60697=>X"00",
60698=>X"00",
60699=>X"00",
60700=>X"00",
60701=>X"00",
60702=>X"00",
60703=>X"00",
60704=>X"00",
60705=>X"00",
60706=>X"00",
60707=>X"00",
60708=>X"00",
60709=>X"00",
60710=>X"00",
60711=>X"00",
60712=>X"00",
60713=>X"00",
60714=>X"00",
60715=>X"00",
60716=>X"00",
60717=>X"00",
60718=>X"00",
60719=>X"00",
60720=>X"00",
60721=>X"00",
60722=>X"00",
60723=>X"00",
60724=>X"00",
60725=>X"00",
60726=>X"00",
60727=>X"00",
60728=>X"00",
60729=>X"00",
60730=>X"00",
60731=>X"00",
60732=>X"00",
60733=>X"00",
60734=>X"00",
60735=>X"00",
60736=>X"00",
60737=>X"00",
60738=>X"00",
60739=>X"00",
60740=>X"00",
60741=>X"00",
60742=>X"00",
60743=>X"00",
60744=>X"00",
60745=>X"00",
60746=>X"00",
60747=>X"00",
60748=>X"00",
60749=>X"00",
60750=>X"00",
60751=>X"00",
60752=>X"00",
60753=>X"00",
60754=>X"00",
60755=>X"00",
60756=>X"00",
60757=>X"00",
60758=>X"00",
60759=>X"00",
60760=>X"00",
60761=>X"00",
60762=>X"00",
60763=>X"00",
60764=>X"00",
60765=>X"00",
60766=>X"00",
60767=>X"00",
60768=>X"00",
60769=>X"00",
60770=>X"00",
60771=>X"00",
60772=>X"00",
60773=>X"00",
60774=>X"00",
60775=>X"00",
60776=>X"00",
60777=>X"00",
60778=>X"00",
60779=>X"00",
60780=>X"00",
60781=>X"00",
60782=>X"00",
60783=>X"00",
60784=>X"00",
60785=>X"00",
60786=>X"00",
60787=>X"00",
60788=>X"00",
60789=>X"00",
60790=>X"00",
60791=>X"00",
60792=>X"00",
60793=>X"00",
60794=>X"00",
60795=>X"00",
60796=>X"00",
60797=>X"00",
60798=>X"00",
60799=>X"00",
60800=>X"00",
60801=>X"00",
60802=>X"00",
60803=>X"00",
60804=>X"00",
60805=>X"00",
60806=>X"00",
60807=>X"00",
60808=>X"00",
60809=>X"00",
60810=>X"00",
60811=>X"00",
60812=>X"00",
60813=>X"00",
60814=>X"00",
60815=>X"00",
60816=>X"00",
60817=>X"00",
60818=>X"00",
60819=>X"00",
60820=>X"00",
60821=>X"00",
60822=>X"00",
60823=>X"00",
60824=>X"00",
60825=>X"00",
60826=>X"00",
60827=>X"00",
60828=>X"00",
60829=>X"00",
60830=>X"00",
60831=>X"00",
60832=>X"00",
60833=>X"00",
60834=>X"00",
60835=>X"00",
60836=>X"00",
60837=>X"00",
60838=>X"00",
60839=>X"00",
60840=>X"00",
60841=>X"00",
60842=>X"00",
60843=>X"00",
60844=>X"00",
60845=>X"00",
60846=>X"00",
60847=>X"00",
60848=>X"00",
60849=>X"00",
60850=>X"00",
60851=>X"00",
60852=>X"00",
60853=>X"00",
60854=>X"00",
60855=>X"00",
60856=>X"00",
60857=>X"00",
60858=>X"00",
60859=>X"00",
60860=>X"00",
60861=>X"00",
60862=>X"00",
60863=>X"00",
60864=>X"00",
60865=>X"00",
60866=>X"00",
60867=>X"00",
60868=>X"00",
60869=>X"00",
60870=>X"00",
60871=>X"00",
60872=>X"00",
60873=>X"00",
60874=>X"00",
60875=>X"00",
60876=>X"00",
60877=>X"00",
60878=>X"00",
60879=>X"00",
60880=>X"00",
60881=>X"00",
60882=>X"00",
60883=>X"00",
60884=>X"00",
60885=>X"00",
60886=>X"00",
60887=>X"00",
60888=>X"00",
60889=>X"00",
60890=>X"00",
60891=>X"00",
60892=>X"00",
60893=>X"00",
60894=>X"00",
60895=>X"00",
60896=>X"00",
60897=>X"00",
60898=>X"00",
60899=>X"00",
60900=>X"00",
60901=>X"00",
60902=>X"00",
60903=>X"00",
60904=>X"00",
60905=>X"00",
60906=>X"00",
60907=>X"00",
60908=>X"00",
60909=>X"00",
60910=>X"00",
60911=>X"00",
60912=>X"00",
60913=>X"00",
60914=>X"00",
60915=>X"00",
60916=>X"00",
60917=>X"00",
60918=>X"00",
60919=>X"00",
60920=>X"00",
60921=>X"00",
60922=>X"00",
60923=>X"00",
60924=>X"00",
60925=>X"00",
60926=>X"00",
60927=>X"00",
60928=>X"00",
60929=>X"00",
60930=>X"00",
60931=>X"00",
60932=>X"00",
60933=>X"00",
60934=>X"00",
60935=>X"00",
60936=>X"00",
60937=>X"00",
60938=>X"00",
60939=>X"00",
60940=>X"00",
60941=>X"00",
60942=>X"00",
60943=>X"00",
60944=>X"00",
60945=>X"00",
60946=>X"00",
60947=>X"00",
60948=>X"00",
60949=>X"00",
60950=>X"00",
60951=>X"00",
60952=>X"00",
60953=>X"00",
60954=>X"00",
60955=>X"00",
60956=>X"00",
60957=>X"00",
60958=>X"00",
60959=>X"00",
60960=>X"00",
60961=>X"00",
60962=>X"00",
60963=>X"00",
60964=>X"00",
60965=>X"00",
60966=>X"00",
60967=>X"00",
60968=>X"00",
60969=>X"00",
60970=>X"00",
60971=>X"00",
60972=>X"00",
60973=>X"00",
60974=>X"00",
60975=>X"00",
60976=>X"00",
60977=>X"00",
60978=>X"00",
60979=>X"00",
60980=>X"00",
60981=>X"00",
60982=>X"00",
60983=>X"00",
60984=>X"00",
60985=>X"00",
60986=>X"00",
60987=>X"00",
60988=>X"00",
60989=>X"00",
60990=>X"00",
60991=>X"00",
60992=>X"00",
60993=>X"00",
60994=>X"00",
60995=>X"00",
60996=>X"00",
60997=>X"00",
60998=>X"00",
60999=>X"00",
61000=>X"00",
61001=>X"00",
61002=>X"00",
61003=>X"00",
61004=>X"00",
61005=>X"00",
61006=>X"00",
61007=>X"00",
61008=>X"00",
61009=>X"00",
61010=>X"00",
61011=>X"00",
61012=>X"00",
61013=>X"00",
61014=>X"00",
61015=>X"00",
61016=>X"00",
61017=>X"00",
61018=>X"00",
61019=>X"00",
61020=>X"00",
61021=>X"00",
61022=>X"00",
61023=>X"00",
61024=>X"00",
61025=>X"00",
61026=>X"00",
61027=>X"00",
61028=>X"00",
61029=>X"00",
61030=>X"00",
61031=>X"00",
61032=>X"00",
61033=>X"00",
61034=>X"00",
61035=>X"00",
61036=>X"00",
61037=>X"00",
61038=>X"00",
61039=>X"00",
61040=>X"00",
61041=>X"00",
61042=>X"00",
61043=>X"00",
61044=>X"00",
61045=>X"00",
61046=>X"00",
61047=>X"00",
61048=>X"00",
61049=>X"00",
61050=>X"00",
61051=>X"00",
61052=>X"00",
61053=>X"00",
61054=>X"00",
61055=>X"00",
61056=>X"00",
61057=>X"00",
61058=>X"00",
61059=>X"00",
61060=>X"00",
61061=>X"00",
61062=>X"00",
61063=>X"00",
61064=>X"00",
61065=>X"00",
61066=>X"00",
61067=>X"00",
61068=>X"00",
61069=>X"00",
61070=>X"00",
61071=>X"00",
61072=>X"00",
61073=>X"00",
61074=>X"00",
61075=>X"00",
61076=>X"00",
61077=>X"00",
61078=>X"00",
61079=>X"00",
61080=>X"00",
61081=>X"00",
61082=>X"00",
61083=>X"00",
61084=>X"00",
61085=>X"00",
61086=>X"00",
61087=>X"00",
61088=>X"00",
61089=>X"00",
61090=>X"00",
61091=>X"00",
61092=>X"00",
61093=>X"00",
61094=>X"00",
61095=>X"00",
61096=>X"00",
61097=>X"00",
61098=>X"00",
61099=>X"00",
61100=>X"00",
61101=>X"00",
61102=>X"00",
61103=>X"00",
61104=>X"00",
61105=>X"00",
61106=>X"00",
61107=>X"00",
61108=>X"00",
61109=>X"00",
61110=>X"00",
61111=>X"00",
61112=>X"00",
61113=>X"00",
61114=>X"00",
61115=>X"00",
61116=>X"00",
61117=>X"00",
61118=>X"00",
61119=>X"00",
61120=>X"00",
61121=>X"00",
61122=>X"00",
61123=>X"00",
61124=>X"00",
61125=>X"00",
61126=>X"00",
61127=>X"00",
61128=>X"00",
61129=>X"00",
61130=>X"00",
61131=>X"00",
61132=>X"00",
61133=>X"00",
61134=>X"00",
61135=>X"00",
61136=>X"00",
61137=>X"00",
61138=>X"00",
61139=>X"00",
61140=>X"00",
61141=>X"00",
61142=>X"00",
61143=>X"00",
61144=>X"00",
61145=>X"00",
61146=>X"00",
61147=>X"00",
61148=>X"00",
61149=>X"00",
61150=>X"00",
61151=>X"00",
61152=>X"00",
61153=>X"00",
61154=>X"00",
61155=>X"00",
61156=>X"00",
61157=>X"00",
61158=>X"00",
61159=>X"00",
61160=>X"00",
61161=>X"00",
61162=>X"00",
61163=>X"00",
61164=>X"00",
61165=>X"00",
61166=>X"00",
61167=>X"00",
61168=>X"00",
61169=>X"00",
61170=>X"00",
61171=>X"00",
61172=>X"00",
61173=>X"00",
61174=>X"00",
61175=>X"00",
61176=>X"00",
61177=>X"00",
61178=>X"00",
61179=>X"00",
61180=>X"00",
61181=>X"00",
61182=>X"00",
61183=>X"00",
61184=>X"00",
61185=>X"00",
61186=>X"00",
61187=>X"00",
61188=>X"00",
61189=>X"00",
61190=>X"00",
61191=>X"00",
61192=>X"00",
61193=>X"00",
61194=>X"00",
61195=>X"00",
61196=>X"00",
61197=>X"00",
61198=>X"00",
61199=>X"00",
61200=>X"00",
61201=>X"00",
61202=>X"00",
61203=>X"00",
61204=>X"00",
61205=>X"00",
61206=>X"00",
61207=>X"00",
61208=>X"00",
61209=>X"00",
61210=>X"00",
61211=>X"00",
61212=>X"00",
61213=>X"00",
61214=>X"00",
61215=>X"00",
61216=>X"00",
61217=>X"00",
61218=>X"00",
61219=>X"00",
61220=>X"00",
61221=>X"00",
61222=>X"00",
61223=>X"00",
61224=>X"00",
61225=>X"00",
61226=>X"00",
61227=>X"00",
61228=>X"00",
61229=>X"00",
61230=>X"00",
61231=>X"00",
61232=>X"00",
61233=>X"00",
61234=>X"00",
61235=>X"00",
61236=>X"00",
61237=>X"00",
61238=>X"00",
61239=>X"00",
61240=>X"00",
61241=>X"00",
61242=>X"00",
61243=>X"00",
61244=>X"00",
61245=>X"00",
61246=>X"00",
61247=>X"00",
61248=>X"00",
61249=>X"00",
61250=>X"00",
61251=>X"00",
61252=>X"00",
61253=>X"00",
61254=>X"00",
61255=>X"00",
61256=>X"00",
61257=>X"00",
61258=>X"00",
61259=>X"00",
61260=>X"00",
61261=>X"00",
61262=>X"00",
61263=>X"00",
61264=>X"00",
61265=>X"00",
61266=>X"00",
61267=>X"00",
61268=>X"00",
61269=>X"00",
61270=>X"00",
61271=>X"00",
61272=>X"00",
61273=>X"00",
61274=>X"00",
61275=>X"00",
61276=>X"00",
61277=>X"00",
61278=>X"00",
61279=>X"00",
61280=>X"00",
61281=>X"00",
61282=>X"00",
61283=>X"00",
61284=>X"00",
61285=>X"00",
61286=>X"00",
61287=>X"00",
61288=>X"00",
61289=>X"00",
61290=>X"00",
61291=>X"00",
61292=>X"00",
61293=>X"00",
61294=>X"00",
61295=>X"00",
61296=>X"00",
61297=>X"00",
61298=>X"00",
61299=>X"00",
61300=>X"00",
61301=>X"00",
61302=>X"00",
61303=>X"00",
61304=>X"00",
61305=>X"00",
61306=>X"00",
61307=>X"00",
61308=>X"00",
61309=>X"00",
61310=>X"00",
61311=>X"00",
61312=>X"00",
61313=>X"00",
61314=>X"00",
61315=>X"00",
61316=>X"00",
61317=>X"00",
61318=>X"00",
61319=>X"00",
61320=>X"00",
61321=>X"00",
61322=>X"00",
61323=>X"00",
61324=>X"00",
61325=>X"00",
61326=>X"00",
61327=>X"00",
61328=>X"00",
61329=>X"00",
61330=>X"00",
61331=>X"00",
61332=>X"00",
61333=>X"00",
61334=>X"00",
61335=>X"00",
61336=>X"00",
61337=>X"00",
61338=>X"00",
61339=>X"00",
61340=>X"00",
61341=>X"00",
61342=>X"00",
61343=>X"00",
61344=>X"00",
61345=>X"00",
61346=>X"00",
61347=>X"00",
61348=>X"00",
61349=>X"00",
61350=>X"00",
61351=>X"00",
61352=>X"00",
61353=>X"00",
61354=>X"00",
61355=>X"00",
61356=>X"00",
61357=>X"00",
61358=>X"00",
61359=>X"00",
61360=>X"00",
61361=>X"00",
61362=>X"00",
61363=>X"00",
61364=>X"00",
61365=>X"00",
61366=>X"00",
61367=>X"00",
61368=>X"00",
61369=>X"00",
61370=>X"00",
61371=>X"00",
61372=>X"00",
61373=>X"00",
61374=>X"00",
61375=>X"00",
61376=>X"00",
61377=>X"00",
61378=>X"00",
61379=>X"00",
61380=>X"00",
61381=>X"00",
61382=>X"00",
61383=>X"00",
61384=>X"00",
61385=>X"00",
61386=>X"00",
61387=>X"00",
61388=>X"00",
61389=>X"00",
61390=>X"00",
61391=>X"00",
61392=>X"00",
61393=>X"00",
61394=>X"00",
61395=>X"00",
61396=>X"00",
61397=>X"00",
61398=>X"00",
61399=>X"00",
61400=>X"00",
61401=>X"00",
61402=>X"00",
61403=>X"00",
61404=>X"00",
61405=>X"00",
61406=>X"00",
61407=>X"00",
61408=>X"00",
61409=>X"00",
61410=>X"00",
61411=>X"00",
61412=>X"00",
61413=>X"00",
61414=>X"00",
61415=>X"00",
61416=>X"00",
61417=>X"00",
61418=>X"00",
61419=>X"00",
61420=>X"00",
61421=>X"00",
61422=>X"00",
61423=>X"00",
61424=>X"00",
61425=>X"00",
61426=>X"00",
61427=>X"00",
61428=>X"00",
61429=>X"00",
61430=>X"00",
61431=>X"00",
61432=>X"00",
61433=>X"00",
61434=>X"00",
61435=>X"00",
61436=>X"00",
61437=>X"00",
61438=>X"00",
61439=>X"00",
61440=>X"00",
61441=>X"00",
61442=>X"00",
61443=>X"00",
61444=>X"00",
61445=>X"00",
61446=>X"00",
61447=>X"00",
61448=>X"00",
61449=>X"00",
61450=>X"00",
61451=>X"00",
61452=>X"00",
61453=>X"00",
61454=>X"00",
61455=>X"00",
61456=>X"00",
61457=>X"00",
61458=>X"00",
61459=>X"00",
61460=>X"00",
61461=>X"00",
61462=>X"00",
61463=>X"00",
61464=>X"00",
61465=>X"00",
61466=>X"00",
61467=>X"00",
61468=>X"00",
61469=>X"00",
61470=>X"00",
61471=>X"00",
61472=>X"00",
61473=>X"00",
61474=>X"00",
61475=>X"00",
61476=>X"00",
61477=>X"00",
61478=>X"00",
61479=>X"00",
61480=>X"00",
61481=>X"00",
61482=>X"00",
61483=>X"00",
61484=>X"00",
61485=>X"00",
61486=>X"00",
61487=>X"00",
61488=>X"00",
61489=>X"00",
61490=>X"00",
61491=>X"00",
61492=>X"00",
61493=>X"00",
61494=>X"00",
61495=>X"00",
61496=>X"00",
61497=>X"00",
61498=>X"00",
61499=>X"00",
61500=>X"00",
61501=>X"00",
61502=>X"00",
61503=>X"00",
61504=>X"00",
61505=>X"00",
61506=>X"00",
61507=>X"00",
61508=>X"00",
61509=>X"00",
61510=>X"00",
61511=>X"00",
61512=>X"00",
61513=>X"00",
61514=>X"00",
61515=>X"00",
61516=>X"00",
61517=>X"00",
61518=>X"00",
61519=>X"00",
61520=>X"00",
61521=>X"00",
61522=>X"00",
61523=>X"00",
61524=>X"00",
61525=>X"00",
61526=>X"00",
61527=>X"00",
61528=>X"00",
61529=>X"00",
61530=>X"00",
61531=>X"00",
61532=>X"00",
61533=>X"00",
61534=>X"00",
61535=>X"00",
61536=>X"00",
61537=>X"00",
61538=>X"00",
61539=>X"00",
61540=>X"00",
61541=>X"00",
61542=>X"00",
61543=>X"00",
61544=>X"00",
61545=>X"00",
61546=>X"00",
61547=>X"00",
61548=>X"00",
61549=>X"00",
61550=>X"00",
61551=>X"00",
61552=>X"00",
61553=>X"00",
61554=>X"00",
61555=>X"00",
61556=>X"00",
61557=>X"00",
61558=>X"00",
61559=>X"00",
61560=>X"00",
61561=>X"00",
61562=>X"00",
61563=>X"00",
61564=>X"00",
61565=>X"00",
61566=>X"00",
61567=>X"00",
61568=>X"00",
61569=>X"00",
61570=>X"00",
61571=>X"00",
61572=>X"00",
61573=>X"00",
61574=>X"00",
61575=>X"00",
61576=>X"00",
61577=>X"00",
61578=>X"00",
61579=>X"00",
61580=>X"00",
61581=>X"00",
61582=>X"00",
61583=>X"00",
61584=>X"00",
61585=>X"00",
61586=>X"00",
61587=>X"00",
61588=>X"00",
61589=>X"00",
61590=>X"00",
61591=>X"00",
61592=>X"00",
61593=>X"00",
61594=>X"00",
61595=>X"00",
61596=>X"00",
61597=>X"00",
61598=>X"00",
61599=>X"00",
61600=>X"00",
61601=>X"00",
61602=>X"00",
61603=>X"00",
61604=>X"00",
61605=>X"00",
61606=>X"00",
61607=>X"00",
61608=>X"00",
61609=>X"00",
61610=>X"00",
61611=>X"00",
61612=>X"00",
61613=>X"00",
61614=>X"00",
61615=>X"00",
61616=>X"00",
61617=>X"00",
61618=>X"00",
61619=>X"00",
61620=>X"00",
61621=>X"00",
61622=>X"00",
61623=>X"00",
61624=>X"00",
61625=>X"00",
61626=>X"00",
61627=>X"00",
61628=>X"00",
61629=>X"00",
61630=>X"00",
61631=>X"00",
61632=>X"00",
61633=>X"00",
61634=>X"00",
61635=>X"00",
61636=>X"00",
61637=>X"00",
61638=>X"00",
61639=>X"00",
61640=>X"00",
61641=>X"00",
61642=>X"00",
61643=>X"00",
61644=>X"00",
61645=>X"00",
61646=>X"00",
61647=>X"00",
61648=>X"00",
61649=>X"00",
61650=>X"00",
61651=>X"00",
61652=>X"00",
61653=>X"00",
61654=>X"00",
61655=>X"00",
61656=>X"00",
61657=>X"00",
61658=>X"00",
61659=>X"00",
61660=>X"00",
61661=>X"00",
61662=>X"00",
61663=>X"00",
61664=>X"00",
61665=>X"00",
61666=>X"00",
61667=>X"00",
61668=>X"00",
61669=>X"00",
61670=>X"00",
61671=>X"00",
61672=>X"00",
61673=>X"00",
61674=>X"00",
61675=>X"00",
61676=>X"00",
61677=>X"00",
61678=>X"00",
61679=>X"00",
61680=>X"00",
61681=>X"00",
61682=>X"00",
61683=>X"00",
61684=>X"00",
61685=>X"00",
61686=>X"00",
61687=>X"00",
61688=>X"00",
61689=>X"00",
61690=>X"00",
61691=>X"00",
61692=>X"00",
61693=>X"00",
61694=>X"00",
61695=>X"00",
61696=>X"00",
61697=>X"00",
61698=>X"00",
61699=>X"00",
61700=>X"00",
61701=>X"00",
61702=>X"00",
61703=>X"00",
61704=>X"00",
61705=>X"00",
61706=>X"00",
61707=>X"00",
61708=>X"00",
61709=>X"00",
61710=>X"00",
61711=>X"00",
61712=>X"00",
61713=>X"00",
61714=>X"00",
61715=>X"00",
61716=>X"00",
61717=>X"00",
61718=>X"00",
61719=>X"00",
61720=>X"00",
61721=>X"00",
61722=>X"00",
61723=>X"00",
61724=>X"00",
61725=>X"00",
61726=>X"00",
61727=>X"00",
61728=>X"00",
61729=>X"00",
61730=>X"00",
61731=>X"00",
61732=>X"00",
61733=>X"00",
61734=>X"00",
61735=>X"00",
61736=>X"00",
61737=>X"00",
61738=>X"00",
61739=>X"00",
61740=>X"00",
61741=>X"00",
61742=>X"00",
61743=>X"00",
61744=>X"00",
61745=>X"00",
61746=>X"00",
61747=>X"00",
61748=>X"00",
61749=>X"00",
61750=>X"00",
61751=>X"00",
61752=>X"00",
61753=>X"00",
61754=>X"00",
61755=>X"00",
61756=>X"00",
61757=>X"00",
61758=>X"00",
61759=>X"00",
61760=>X"00",
61761=>X"00",
61762=>X"00",
61763=>X"00",
61764=>X"00",
61765=>X"00",
61766=>X"00",
61767=>X"00",
61768=>X"00",
61769=>X"00",
61770=>X"00",
61771=>X"00",
61772=>X"00",
61773=>X"00",
61774=>X"00",
61775=>X"00",
61776=>X"00",
61777=>X"00",
61778=>X"00",
61779=>X"00",
61780=>X"00",
61781=>X"00",
61782=>X"00",
61783=>X"00",
61784=>X"00",
61785=>X"00",
61786=>X"00",
61787=>X"00",
61788=>X"00",
61789=>X"00",
61790=>X"00",
61791=>X"00",
61792=>X"00",
61793=>X"00",
61794=>X"00",
61795=>X"00",
61796=>X"00",
61797=>X"00",
61798=>X"00",
61799=>X"00",
61800=>X"00",
61801=>X"00",
61802=>X"00",
61803=>X"00",
61804=>X"00",
61805=>X"00",
61806=>X"00",
61807=>X"00",
61808=>X"00",
61809=>X"00",
61810=>X"00",
61811=>X"00",
61812=>X"00",
61813=>X"00",
61814=>X"00",
61815=>X"00",
61816=>X"00",
61817=>X"00",
61818=>X"00",
61819=>X"00",
61820=>X"00",
61821=>X"00",
61822=>X"00",
61823=>X"00",
61824=>X"00",
61825=>X"00",
61826=>X"00",
61827=>X"00",
61828=>X"00",
61829=>X"00",
61830=>X"00",
61831=>X"00",
61832=>X"00",
61833=>X"00",
61834=>X"00",
61835=>X"00",
61836=>X"00",
61837=>X"00",
61838=>X"00",
61839=>X"00",
61840=>X"00",
61841=>X"00",
61842=>X"00",
61843=>X"00",
61844=>X"00",
61845=>X"00",
61846=>X"00",
61847=>X"00",
61848=>X"00",
61849=>X"00",
61850=>X"00",
61851=>X"00",
61852=>X"00",
61853=>X"00",
61854=>X"00",
61855=>X"00",
61856=>X"00",
61857=>X"00",
61858=>X"00",
61859=>X"00",
61860=>X"00",
61861=>X"00",
61862=>X"00",
61863=>X"00",
61864=>X"00",
61865=>X"00",
61866=>X"00",
61867=>X"00",
61868=>X"00",
61869=>X"00",
61870=>X"00",
61871=>X"00",
61872=>X"00",
61873=>X"00",
61874=>X"00",
61875=>X"00",
61876=>X"00",
61877=>X"00",
61878=>X"00",
61879=>X"00",
61880=>X"00",
61881=>X"00",
61882=>X"00",
61883=>X"00",
61884=>X"00",
61885=>X"00",
61886=>X"00",
61887=>X"00",
61888=>X"00",
61889=>X"00",
61890=>X"00",
61891=>X"00",
61892=>X"00",
61893=>X"00",
61894=>X"00",
61895=>X"00",
61896=>X"00",
61897=>X"00",
61898=>X"00",
61899=>X"00",
61900=>X"00",
61901=>X"00",
61902=>X"00",
61903=>X"00",
61904=>X"00",
61905=>X"00",
61906=>X"00",
61907=>X"00",
61908=>X"00",
61909=>X"00",
61910=>X"00",
61911=>X"00",
61912=>X"00",
61913=>X"00",
61914=>X"00",
61915=>X"00",
61916=>X"00",
61917=>X"00",
61918=>X"00",
61919=>X"00",
61920=>X"00",
61921=>X"00",
61922=>X"00",
61923=>X"00",
61924=>X"00",
61925=>X"00",
61926=>X"00",
61927=>X"00",
61928=>X"00",
61929=>X"00",
61930=>X"00",
61931=>X"00",
61932=>X"00",
61933=>X"00",
61934=>X"00",
61935=>X"00",
61936=>X"00",
61937=>X"00",
61938=>X"00",
61939=>X"00",
61940=>X"00",
61941=>X"00",
61942=>X"00",
61943=>X"00",
61944=>X"00",
61945=>X"00",
61946=>X"00",
61947=>X"00",
61948=>X"00",
61949=>X"00",
61950=>X"00",
61951=>X"00",
61952=>X"00",
61953=>X"00",
61954=>X"00",
61955=>X"00",
61956=>X"00",
61957=>X"00",
61958=>X"00",
61959=>X"00",
61960=>X"00",
61961=>X"00",
61962=>X"00",
61963=>X"00",
61964=>X"00",
61965=>X"00",
61966=>X"00",
61967=>X"00",
61968=>X"00",
61969=>X"00",
61970=>X"00",
61971=>X"00",
61972=>X"00",
61973=>X"00",
61974=>X"00",
61975=>X"00",
61976=>X"00",
61977=>X"00",
61978=>X"00",
61979=>X"00",
61980=>X"00",
61981=>X"00",
61982=>X"00",
61983=>X"00",
61984=>X"00",
61985=>X"00",
61986=>X"00",
61987=>X"00",
61988=>X"00",
61989=>X"00",
61990=>X"00",
61991=>X"00",
61992=>X"00",
61993=>X"00",
61994=>X"00",
61995=>X"00",
61996=>X"00",
61997=>X"00",
61998=>X"00",
61999=>X"00",
62000=>X"00",
62001=>X"00",
62002=>X"00",
62003=>X"00",
62004=>X"00",
62005=>X"00",
62006=>X"00",
62007=>X"00",
62008=>X"00",
62009=>X"00",
62010=>X"00",
62011=>X"00",
62012=>X"00",
62013=>X"00",
62014=>X"00",
62015=>X"00",
62016=>X"00",
62017=>X"00",
62018=>X"00",
62019=>X"00",
62020=>X"00",
62021=>X"00",
62022=>X"00",
62023=>X"00",
62024=>X"00",
62025=>X"00",
62026=>X"00",
62027=>X"00",
62028=>X"00",
62029=>X"00",
62030=>X"00",
62031=>X"00",
62032=>X"00",
62033=>X"00",
62034=>X"00",
62035=>X"00",
62036=>X"00",
62037=>X"00",
62038=>X"00",
62039=>X"00",
62040=>X"00",
62041=>X"00",
62042=>X"00",
62043=>X"00",
62044=>X"00",
62045=>X"00",
62046=>X"00",
62047=>X"00",
62048=>X"00",
62049=>X"00",
62050=>X"00",
62051=>X"00",
62052=>X"00",
62053=>X"00",
62054=>X"00",
62055=>X"00",
62056=>X"00",
62057=>X"00",
62058=>X"00",
62059=>X"00",
62060=>X"00",
62061=>X"00",
62062=>X"00",
62063=>X"00",
62064=>X"00",
62065=>X"00",
62066=>X"00",
62067=>X"00",
62068=>X"00",
62069=>X"00",
62070=>X"00",
62071=>X"00",
62072=>X"00",
62073=>X"00",
62074=>X"00",
62075=>X"00",
62076=>X"00",
62077=>X"00",
62078=>X"00",
62079=>X"00",
62080=>X"00",
62081=>X"00",
62082=>X"00",
62083=>X"00",
62084=>X"00",
62085=>X"00",
62086=>X"00",
62087=>X"00",
62088=>X"00",
62089=>X"00",
62090=>X"00",
62091=>X"00",
62092=>X"00",
62093=>X"00",
62094=>X"00",
62095=>X"00",
62096=>X"00",
62097=>X"00",
62098=>X"00",
62099=>X"00",
62100=>X"00",
62101=>X"00",
62102=>X"00",
62103=>X"00",
62104=>X"00",
62105=>X"00",
62106=>X"00",
62107=>X"00",
62108=>X"00",
62109=>X"00",
62110=>X"00",
62111=>X"00",
62112=>X"00",
62113=>X"00",
62114=>X"00",
62115=>X"00",
62116=>X"00",
62117=>X"00",
62118=>X"00",
62119=>X"00",
62120=>X"00",
62121=>X"00",
62122=>X"00",
62123=>X"00",
62124=>X"00",
62125=>X"00",
62126=>X"00",
62127=>X"00",
62128=>X"00",
62129=>X"00",
62130=>X"00",
62131=>X"00",
62132=>X"00",
62133=>X"00",
62134=>X"00",
62135=>X"00",
62136=>X"00",
62137=>X"00",
62138=>X"00",
62139=>X"00",
62140=>X"00",
62141=>X"00",
62142=>X"00",
62143=>X"00",
62144=>X"00",
62145=>X"00",
62146=>X"00",
62147=>X"00",
62148=>X"00",
62149=>X"00",
62150=>X"00",
62151=>X"00",
62152=>X"00",
62153=>X"00",
62154=>X"00",
62155=>X"00",
62156=>X"00",
62157=>X"00",
62158=>X"00",
62159=>X"00",
62160=>X"00",
62161=>X"00",
62162=>X"00",
62163=>X"00",
62164=>X"00",
62165=>X"00",
62166=>X"00",
62167=>X"00",
62168=>X"00",
62169=>X"00",
62170=>X"00",
62171=>X"00",
62172=>X"00",
62173=>X"00",
62174=>X"00",
62175=>X"00",
62176=>X"00",
62177=>X"00",
62178=>X"00",
62179=>X"00",
62180=>X"00",
62181=>X"00",
62182=>X"00",
62183=>X"00",
62184=>X"00",
62185=>X"00",
62186=>X"00",
62187=>X"00",
62188=>X"00",
62189=>X"00",
62190=>X"00",
62191=>X"00",
62192=>X"00",
62193=>X"00",
62194=>X"00",
62195=>X"00",
62196=>X"00",
62197=>X"00",
62198=>X"00",
62199=>X"00",
62200=>X"00",
62201=>X"00",
62202=>X"00",
62203=>X"00",
62204=>X"00",
62205=>X"00",
62206=>X"00",
62207=>X"00",
62208=>X"00",
62209=>X"00",
62210=>X"00",
62211=>X"00",
62212=>X"00",
62213=>X"00",
62214=>X"00",
62215=>X"00",
62216=>X"00",
62217=>X"00",
62218=>X"00",
62219=>X"00",
62220=>X"00",
62221=>X"00",
62222=>X"00",
62223=>X"00",
62224=>X"00",
62225=>X"00",
62226=>X"00",
62227=>X"00",
62228=>X"00",
62229=>X"00",
62230=>X"00",
62231=>X"00",
62232=>X"00",
62233=>X"00",
62234=>X"00",
62235=>X"00",
62236=>X"00",
62237=>X"00",
62238=>X"00",
62239=>X"00",
62240=>X"00",
62241=>X"00",
62242=>X"00",
62243=>X"00",
62244=>X"00",
62245=>X"00",
62246=>X"00",
62247=>X"00",
62248=>X"00",
62249=>X"00",
62250=>X"00",
62251=>X"00",
62252=>X"00",
62253=>X"00",
62254=>X"00",
62255=>X"00",
62256=>X"00",
62257=>X"00",
62258=>X"00",
62259=>X"00",
62260=>X"00",
62261=>X"00",
62262=>X"00",
62263=>X"00",
62264=>X"00",
62265=>X"00",
62266=>X"00",
62267=>X"00",
62268=>X"00",
62269=>X"00",
62270=>X"00",
62271=>X"00",
62272=>X"00",
62273=>X"00",
62274=>X"00",
62275=>X"00",
62276=>X"00",
62277=>X"00",
62278=>X"00",
62279=>X"00",
62280=>X"00",
62281=>X"00",
62282=>X"00",
62283=>X"00",
62284=>X"00",
62285=>X"00",
62286=>X"00",
62287=>X"00",
62288=>X"00",
62289=>X"00",
62290=>X"00",
62291=>X"00",
62292=>X"00",
62293=>X"00",
62294=>X"00",
62295=>X"00",
62296=>X"00",
62297=>X"00",
62298=>X"00",
62299=>X"00",
62300=>X"00",
62301=>X"00",
62302=>X"00",
62303=>X"00",
62304=>X"00",
62305=>X"00",
62306=>X"00",
62307=>X"00",
62308=>X"00",
62309=>X"00",
62310=>X"00",
62311=>X"00",
62312=>X"00",
62313=>X"00",
62314=>X"00",
62315=>X"00",
62316=>X"00",
62317=>X"00",
62318=>X"00",
62319=>X"00",
62320=>X"00",
62321=>X"00",
62322=>X"00",
62323=>X"00",
62324=>X"00",
62325=>X"00",
62326=>X"00",
62327=>X"00",
62328=>X"00",
62329=>X"00",
62330=>X"00",
62331=>X"00",
62332=>X"00",
62333=>X"00",
62334=>X"00",
62335=>X"00",
62336=>X"00",
62337=>X"00",
62338=>X"00",
62339=>X"00",
62340=>X"00",
62341=>X"00",
62342=>X"00",
62343=>X"00",
62344=>X"00",
62345=>X"00",
62346=>X"00",
62347=>X"00",
62348=>X"00",
62349=>X"00",
62350=>X"00",
62351=>X"00",
62352=>X"00",
62353=>X"00",
62354=>X"00",
62355=>X"00",
62356=>X"00",
62357=>X"00",
62358=>X"00",
62359=>X"00",
62360=>X"00",
62361=>X"00",
62362=>X"00",
62363=>X"00",
62364=>X"00",
62365=>X"00",
62366=>X"00",
62367=>X"00",
62368=>X"00",
62369=>X"00",
62370=>X"00",
62371=>X"00",
62372=>X"00",
62373=>X"00",
62374=>X"00",
62375=>X"00",
62376=>X"00",
62377=>X"00",
62378=>X"00",
62379=>X"00",
62380=>X"00",
62381=>X"00",
62382=>X"00",
62383=>X"00",
62384=>X"00",
62385=>X"00",
62386=>X"00",
62387=>X"00",
62388=>X"00",
62389=>X"00",
62390=>X"00",
62391=>X"00",
62392=>X"00",
62393=>X"00",
62394=>X"00",
62395=>X"00",
62396=>X"00",
62397=>X"00",
62398=>X"00",
62399=>X"00",
62400=>X"00",
62401=>X"00",
62402=>X"00",
62403=>X"00",
62404=>X"00",
62405=>X"00",
62406=>X"00",
62407=>X"00",
62408=>X"00",
62409=>X"00",
62410=>X"00",
62411=>X"00",
62412=>X"00",
62413=>X"00",
62414=>X"00",
62415=>X"00",
62416=>X"00",
62417=>X"00",
62418=>X"00",
62419=>X"00",
62420=>X"00",
62421=>X"00",
62422=>X"00",
62423=>X"00",
62424=>X"00",
62425=>X"00",
62426=>X"00",
62427=>X"00",
62428=>X"00",
62429=>X"00",
62430=>X"00",
62431=>X"00",
62432=>X"00",
62433=>X"00",
62434=>X"00",
62435=>X"00",
62436=>X"00",
62437=>X"00",
62438=>X"00",
62439=>X"00",
62440=>X"00",
62441=>X"00",
62442=>X"00",
62443=>X"00",
62444=>X"00",
62445=>X"00",
62446=>X"00",
62447=>X"00",
62448=>X"00",
62449=>X"00",
62450=>X"00",
62451=>X"00",
62452=>X"00",
62453=>X"00",
62454=>X"00",
62455=>X"00",
62456=>X"00",
62457=>X"00",
62458=>X"00",
62459=>X"00",
62460=>X"00",
62461=>X"00",
62462=>X"00",
62463=>X"00",
62464=>X"00",
62465=>X"00",
62466=>X"00",
62467=>X"00",
62468=>X"00",
62469=>X"00",
62470=>X"00",
62471=>X"00",
62472=>X"00",
62473=>X"00",
62474=>X"00",
62475=>X"00",
62476=>X"00",
62477=>X"00",
62478=>X"00",
62479=>X"00",
62480=>X"00",
62481=>X"00",
62482=>X"00",
62483=>X"00",
62484=>X"00",
62485=>X"00",
62486=>X"00",
62487=>X"00",
62488=>X"00",
62489=>X"00",
62490=>X"00",
62491=>X"00",
62492=>X"00",
62493=>X"00",
62494=>X"00",
62495=>X"00",
62496=>X"00",
62497=>X"00",
62498=>X"00",
62499=>X"00",
62500=>X"00",
62501=>X"00",
62502=>X"00",
62503=>X"00",
62504=>X"00",
62505=>X"00",
62506=>X"00",
62507=>X"00",
62508=>X"00",
62509=>X"00",
62510=>X"00",
62511=>X"00",
62512=>X"00",
62513=>X"00",
62514=>X"00",
62515=>X"00",
62516=>X"00",
62517=>X"00",
62518=>X"00",
62519=>X"00",
62520=>X"00",
62521=>X"00",
62522=>X"00",
62523=>X"00",
62524=>X"00",
62525=>X"00",
62526=>X"00",
62527=>X"00",
62528=>X"00",
62529=>X"00",
62530=>X"00",
62531=>X"00",
62532=>X"00",
62533=>X"00",
62534=>X"00",
62535=>X"00",
62536=>X"00",
62537=>X"00",
62538=>X"00",
62539=>X"00",
62540=>X"00",
62541=>X"00",
62542=>X"00",
62543=>X"00",
62544=>X"00",
62545=>X"00",
62546=>X"00",
62547=>X"00",
62548=>X"00",
62549=>X"00",
62550=>X"00",
62551=>X"00",
62552=>X"00",
62553=>X"00",
62554=>X"00",
62555=>X"00",
62556=>X"00",
62557=>X"00",
62558=>X"00",
62559=>X"00",
62560=>X"00",
62561=>X"00",
62562=>X"00",
62563=>X"00",
62564=>X"00",
62565=>X"00",
62566=>X"00",
62567=>X"00",
62568=>X"00",
62569=>X"00",
62570=>X"00",
62571=>X"00",
62572=>X"00",
62573=>X"00",
62574=>X"00",
62575=>X"00",
62576=>X"00",
62577=>X"00",
62578=>X"00",
62579=>X"00",
62580=>X"00",
62581=>X"00",
62582=>X"00",
62583=>X"00",
62584=>X"00",
62585=>X"00",
62586=>X"00",
62587=>X"00",
62588=>X"00",
62589=>X"00",
62590=>X"00",
62591=>X"00",
62592=>X"00",
62593=>X"00",
62594=>X"00",
62595=>X"00",
62596=>X"00",
62597=>X"00",
62598=>X"00",
62599=>X"00",
62600=>X"00",
62601=>X"00",
62602=>X"00",
62603=>X"00",
62604=>X"00",
62605=>X"00",
62606=>X"00",
62607=>X"00",
62608=>X"00",
62609=>X"00",
62610=>X"00",
62611=>X"00",
62612=>X"00",
62613=>X"00",
62614=>X"00",
62615=>X"00",
62616=>X"00",
62617=>X"00",
62618=>X"00",
62619=>X"00",
62620=>X"00",
62621=>X"00",
62622=>X"00",
62623=>X"00",
62624=>X"00",
62625=>X"00",
62626=>X"00",
62627=>X"00",
62628=>X"00",
62629=>X"00",
62630=>X"00",
62631=>X"00",
62632=>X"00",
62633=>X"00",
62634=>X"00",
62635=>X"00",
62636=>X"00",
62637=>X"00",
62638=>X"00",
62639=>X"00",
62640=>X"00",
62641=>X"00",
62642=>X"00",
62643=>X"00",
62644=>X"00",
62645=>X"00",
62646=>X"00",
62647=>X"00",
62648=>X"00",
62649=>X"00",
62650=>X"00",
62651=>X"00",
62652=>X"00",
62653=>X"00",
62654=>X"00",
62655=>X"00",
62656=>X"00",
62657=>X"00",
62658=>X"00",
62659=>X"00",
62660=>X"00",
62661=>X"00",
62662=>X"00",
62663=>X"00",
62664=>X"00",
62665=>X"00",
62666=>X"00",
62667=>X"00",
62668=>X"00",
62669=>X"00",
62670=>X"00",
62671=>X"00",
62672=>X"00",
62673=>X"00",
62674=>X"00",
62675=>X"00",
62676=>X"00",
62677=>X"00",
62678=>X"00",
62679=>X"00",
62680=>X"00",
62681=>X"00",
62682=>X"00",
62683=>X"00",
62684=>X"00",
62685=>X"00",
62686=>X"00",
62687=>X"00",
62688=>X"00",
62689=>X"00",
62690=>X"00",
62691=>X"00",
62692=>X"00",
62693=>X"00",
62694=>X"00",
62695=>X"00",
62696=>X"00",
62697=>X"00",
62698=>X"00",
62699=>X"00",
62700=>X"00",
62701=>X"00",
62702=>X"00",
62703=>X"00",
62704=>X"00",
62705=>X"00",
62706=>X"00",
62707=>X"00",
62708=>X"00",
62709=>X"00",
62710=>X"00",
62711=>X"00",
62712=>X"00",
62713=>X"00",
62714=>X"00",
62715=>X"00",
62716=>X"00",
62717=>X"00",
62718=>X"00",
62719=>X"00",
62720=>X"00",
62721=>X"00",
62722=>X"00",
62723=>X"00",
62724=>X"00",
62725=>X"00",
62726=>X"00",
62727=>X"00",
62728=>X"00",
62729=>X"00",
62730=>X"00",
62731=>X"00",
62732=>X"00",
62733=>X"00",
62734=>X"00",
62735=>X"00",
62736=>X"00",
62737=>X"00",
62738=>X"00",
62739=>X"00",
62740=>X"00",
62741=>X"00",
62742=>X"00",
62743=>X"00",
62744=>X"00",
62745=>X"00",
62746=>X"00",
62747=>X"00",
62748=>X"00",
62749=>X"00",
62750=>X"00",
62751=>X"00",
62752=>X"00",
62753=>X"00",
62754=>X"00",
62755=>X"00",
62756=>X"00",
62757=>X"00",
62758=>X"00",
62759=>X"00",
62760=>X"00",
62761=>X"00",
62762=>X"00",
62763=>X"00",
62764=>X"00",
62765=>X"00",
62766=>X"00",
62767=>X"00",
62768=>X"00",
62769=>X"00",
62770=>X"00",
62771=>X"00",
62772=>X"00",
62773=>X"00",
62774=>X"00",
62775=>X"00",
62776=>X"00",
62777=>X"00",
62778=>X"00",
62779=>X"00",
62780=>X"00",
62781=>X"00",
62782=>X"00",
62783=>X"00",
62784=>X"00",
62785=>X"00",
62786=>X"00",
62787=>X"00",
62788=>X"00",
62789=>X"00",
62790=>X"00",
62791=>X"00",
62792=>X"00",
62793=>X"00",
62794=>X"00",
62795=>X"00",
62796=>X"00",
62797=>X"00",
62798=>X"00",
62799=>X"00",
62800=>X"00",
62801=>X"00",
62802=>X"00",
62803=>X"00",
62804=>X"00",
62805=>X"00",
62806=>X"00",
62807=>X"00",
62808=>X"00",
62809=>X"00",
62810=>X"00",
62811=>X"00",
62812=>X"00",
62813=>X"00",
62814=>X"00",
62815=>X"00",
62816=>X"00",
62817=>X"00",
62818=>X"00",
62819=>X"00",
62820=>X"00",
62821=>X"00",
62822=>X"00",
62823=>X"00",
62824=>X"00",
62825=>X"00",
62826=>X"00",
62827=>X"00",
62828=>X"00",
62829=>X"00",
62830=>X"00",
62831=>X"00",
62832=>X"00",
62833=>X"00",
62834=>X"00",
62835=>X"00",
62836=>X"00",
62837=>X"00",
62838=>X"00",
62839=>X"00",
62840=>X"00",
62841=>X"00",
62842=>X"00",
62843=>X"00",
62844=>X"00",
62845=>X"00",
62846=>X"00",
62847=>X"00",
62848=>X"00",
62849=>X"00",
62850=>X"00",
62851=>X"00",
62852=>X"00",
62853=>X"00",
62854=>X"00",
62855=>X"00",
62856=>X"00",
62857=>X"00",
62858=>X"00",
62859=>X"00",
62860=>X"00",
62861=>X"00",
62862=>X"00",
62863=>X"00",
62864=>X"00",
62865=>X"00",
62866=>X"00",
62867=>X"00",
62868=>X"00",
62869=>X"00",
62870=>X"00",
62871=>X"00",
62872=>X"00",
62873=>X"00",
62874=>X"00",
62875=>X"00",
62876=>X"00",
62877=>X"00",
62878=>X"00",
62879=>X"00",
62880=>X"00",
62881=>X"00",
62882=>X"00",
62883=>X"00",
62884=>X"00",
62885=>X"00",
62886=>X"00",
62887=>X"00",
62888=>X"00",
62889=>X"00",
62890=>X"00",
62891=>X"00",
62892=>X"00",
62893=>X"00",
62894=>X"00",
62895=>X"00",
62896=>X"00",
62897=>X"00",
62898=>X"00",
62899=>X"00",
62900=>X"00",
62901=>X"00",
62902=>X"00",
62903=>X"00",
62904=>X"00",
62905=>X"00",
62906=>X"00",
62907=>X"00",
62908=>X"00",
62909=>X"00",
62910=>X"00",
62911=>X"00",
62912=>X"00",
62913=>X"00",
62914=>X"00",
62915=>X"00",
62916=>X"00",
62917=>X"00",
62918=>X"00",
62919=>X"00",
62920=>X"00",
62921=>X"00",
62922=>X"00",
62923=>X"00",
62924=>X"00",
62925=>X"00",
62926=>X"00",
62927=>X"00",
62928=>X"00",
62929=>X"00",
62930=>X"00",
62931=>X"00",
62932=>X"00",
62933=>X"00",
62934=>X"00",
62935=>X"00",
62936=>X"00",
62937=>X"00",
62938=>X"00",
62939=>X"00",
62940=>X"00",
62941=>X"00",
62942=>X"00",
62943=>X"00",
62944=>X"00",
62945=>X"00",
62946=>X"00",
62947=>X"00",
62948=>X"00",
62949=>X"00",
62950=>X"00",
62951=>X"00",
62952=>X"00",
62953=>X"00",
62954=>X"00",
62955=>X"00",
62956=>X"00",
62957=>X"00",
62958=>X"00",
62959=>X"00",
62960=>X"00",
62961=>X"00",
62962=>X"00",
62963=>X"00",
62964=>X"00",
62965=>X"00",
62966=>X"00",
62967=>X"00",
62968=>X"00",
62969=>X"00",
62970=>X"00",
62971=>X"00",
62972=>X"00",
62973=>X"00",
62974=>X"00",
62975=>X"00",
62976=>X"00",
62977=>X"00",
62978=>X"00",
62979=>X"00",
62980=>X"00",
62981=>X"00",
62982=>X"00",
62983=>X"00",
62984=>X"00",
62985=>X"00",
62986=>X"00",
62987=>X"00",
62988=>X"00",
62989=>X"00",
62990=>X"00",
62991=>X"00",
62992=>X"00",
62993=>X"00",
62994=>X"00",
62995=>X"00",
62996=>X"00",
62997=>X"00",
62998=>X"00",
62999=>X"00",
63000=>X"00",
63001=>X"00",
63002=>X"00",
63003=>X"00",
63004=>X"00",
63005=>X"00",
63006=>X"00",
63007=>X"00",
63008=>X"00",
63009=>X"00",
63010=>X"00",
63011=>X"00",
63012=>X"00",
63013=>X"00",
63014=>X"00",
63015=>X"00",
63016=>X"00",
63017=>X"00",
63018=>X"00",
63019=>X"00",
63020=>X"00",
63021=>X"00",
63022=>X"00",
63023=>X"00",
63024=>X"00",
63025=>X"00",
63026=>X"00",
63027=>X"00",
63028=>X"00",
63029=>X"00",
63030=>X"00",
63031=>X"00",
63032=>X"00",
63033=>X"00",
63034=>X"00",
63035=>X"00",
63036=>X"00",
63037=>X"00",
63038=>X"00",
63039=>X"00",
63040=>X"00",
63041=>X"00",
63042=>X"00",
63043=>X"00",
63044=>X"00",
63045=>X"00",
63046=>X"00",
63047=>X"00",
63048=>X"00",
63049=>X"00",
63050=>X"00",
63051=>X"00",
63052=>X"00",
63053=>X"00",
63054=>X"00",
63055=>X"00",
63056=>X"00",
63057=>X"00",
63058=>X"00",
63059=>X"00",
63060=>X"00",
63061=>X"00",
63062=>X"00",
63063=>X"00",
63064=>X"00",
63065=>X"00",
63066=>X"00",
63067=>X"00",
63068=>X"00",
63069=>X"00",
63070=>X"00",
63071=>X"00",
63072=>X"00",
63073=>X"00",
63074=>X"00",
63075=>X"00",
63076=>X"00",
63077=>X"00",
63078=>X"00",
63079=>X"00",
63080=>X"00",
63081=>X"00",
63082=>X"00",
63083=>X"00",
63084=>X"00",
63085=>X"00",
63086=>X"00",
63087=>X"00",
63088=>X"00",
63089=>X"00",
63090=>X"00",
63091=>X"00",
63092=>X"00",
63093=>X"00",
63094=>X"00",
63095=>X"00",
63096=>X"00",
63097=>X"00",
63098=>X"00",
63099=>X"00",
63100=>X"00",
63101=>X"00",
63102=>X"00",
63103=>X"00",
63104=>X"00",
63105=>X"00",
63106=>X"00",
63107=>X"00",
63108=>X"00",
63109=>X"00",
63110=>X"00",
63111=>X"00",
63112=>X"00",
63113=>X"00",
63114=>X"00",
63115=>X"00",
63116=>X"00",
63117=>X"00",
63118=>X"00",
63119=>X"00",
63120=>X"00",
63121=>X"00",
63122=>X"00",
63123=>X"00",
63124=>X"00",
63125=>X"00",
63126=>X"00",
63127=>X"00",
63128=>X"00",
63129=>X"00",
63130=>X"00",
63131=>X"00",
63132=>X"00",
63133=>X"00",
63134=>X"00",
63135=>X"00",
63136=>X"00",
63137=>X"00",
63138=>X"00",
63139=>X"00",
63140=>X"00",
63141=>X"00",
63142=>X"00",
63143=>X"00",
63144=>X"00",
63145=>X"00",
63146=>X"00",
63147=>X"00",
63148=>X"00",
63149=>X"00",
63150=>X"00",
63151=>X"00",
63152=>X"00",
63153=>X"00",
63154=>X"00",
63155=>X"00",
63156=>X"00",
63157=>X"00",
63158=>X"00",
63159=>X"00",
63160=>X"00",
63161=>X"00",
63162=>X"00",
63163=>X"00",
63164=>X"00",
63165=>X"00",
63166=>X"00",
63167=>X"00",
63168=>X"00",
63169=>X"00",
63170=>X"00",
63171=>X"00",
63172=>X"00",
63173=>X"00",
63174=>X"00",
63175=>X"00",
63176=>X"00",
63177=>X"00",
63178=>X"00",
63179=>X"00",
63180=>X"00",
63181=>X"00",
63182=>X"00",
63183=>X"00",
63184=>X"00",
63185=>X"00",
63186=>X"00",
63187=>X"00",
63188=>X"00",
63189=>X"00",
63190=>X"00",
63191=>X"00",
63192=>X"00",
63193=>X"00",
63194=>X"00",
63195=>X"00",
63196=>X"00",
63197=>X"00",
63198=>X"00",
63199=>X"00",
63200=>X"00",
63201=>X"00",
63202=>X"00",
63203=>X"00",
63204=>X"00",
63205=>X"00",
63206=>X"00",
63207=>X"00",
63208=>X"00",
63209=>X"00",
63210=>X"00",
63211=>X"00",
63212=>X"00",
63213=>X"00",
63214=>X"00",
63215=>X"00",
63216=>X"00",
63217=>X"00",
63218=>X"00",
63219=>X"00",
63220=>X"00",
63221=>X"00",
63222=>X"00",
63223=>X"00",
63224=>X"00",
63225=>X"00",
63226=>X"00",
63227=>X"00",
63228=>X"00",
63229=>X"00",
63230=>X"00",
63231=>X"00",
63232=>X"00",
63233=>X"00",
63234=>X"00",
63235=>X"00",
63236=>X"00",
63237=>X"00",
63238=>X"00",
63239=>X"00",
63240=>X"00",
63241=>X"00",
63242=>X"00",
63243=>X"00",
63244=>X"00",
63245=>X"00",
63246=>X"00",
63247=>X"00",
63248=>X"00",
63249=>X"00",
63250=>X"00",
63251=>X"00",
63252=>X"00",
63253=>X"00",
63254=>X"00",
63255=>X"00",
63256=>X"00",
63257=>X"00",
63258=>X"00",
63259=>X"00",
63260=>X"00",
63261=>X"00",
63262=>X"00",
63263=>X"00",
63264=>X"00",
63265=>X"00",
63266=>X"00",
63267=>X"00",
63268=>X"00",
63269=>X"00",
63270=>X"00",
63271=>X"00",
63272=>X"00",
63273=>X"00",
63274=>X"00",
63275=>X"00",
63276=>X"00",
63277=>X"00",
63278=>X"00",
63279=>X"00",
63280=>X"00",
63281=>X"00",
63282=>X"00",
63283=>X"00",
63284=>X"00",
63285=>X"00",
63286=>X"00",
63287=>X"00",
63288=>X"00",
63289=>X"00",
63290=>X"00",
63291=>X"00",
63292=>X"00",
63293=>X"00",
63294=>X"00",
63295=>X"00",
63296=>X"00",
63297=>X"00",
63298=>X"00",
63299=>X"00",
63300=>X"00",
63301=>X"00",
63302=>X"00",
63303=>X"00",
63304=>X"00",
63305=>X"00",
63306=>X"00",
63307=>X"00",
63308=>X"00",
63309=>X"00",
63310=>X"00",
63311=>X"00",
63312=>X"00",
63313=>X"00",
63314=>X"00",
63315=>X"00",
63316=>X"00",
63317=>X"00",
63318=>X"00",
63319=>X"00",
63320=>X"00",
63321=>X"00",
63322=>X"00",
63323=>X"00",
63324=>X"00",
63325=>X"00",
63326=>X"00",
63327=>X"00",
63328=>X"00",
63329=>X"00",
63330=>X"00",
63331=>X"00",
63332=>X"00",
63333=>X"00",
63334=>X"00",
63335=>X"00",
63336=>X"00",
63337=>X"00",
63338=>X"00",
63339=>X"00",
63340=>X"00",
63341=>X"00",
63342=>X"00",
63343=>X"00",
63344=>X"00",
63345=>X"00",
63346=>X"00",
63347=>X"00",
63348=>X"00",
63349=>X"00",
63350=>X"00",
63351=>X"00",
63352=>X"00",
63353=>X"00",
63354=>X"00",
63355=>X"00",
63356=>X"00",
63357=>X"00",
63358=>X"00",
63359=>X"00",
63360=>X"00",
63361=>X"00",
63362=>X"00",
63363=>X"00",
63364=>X"00",
63365=>X"00",
63366=>X"00",
63367=>X"00",
63368=>X"00",
63369=>X"00",
63370=>X"00",
63371=>X"00",
63372=>X"00",
63373=>X"00",
63374=>X"00",
63375=>X"00",
63376=>X"00",
63377=>X"00",
63378=>X"00",
63379=>X"00",
63380=>X"00",
63381=>X"00",
63382=>X"00",
63383=>X"00",
63384=>X"00",
63385=>X"00",
63386=>X"00",
63387=>X"00",
63388=>X"00",
63389=>X"00",
63390=>X"00",
63391=>X"00",
63392=>X"00",
63393=>X"00",
63394=>X"00",
63395=>X"00",
63396=>X"00",
63397=>X"00",
63398=>X"00",
63399=>X"00",
63400=>X"00",
63401=>X"00",
63402=>X"00",
63403=>X"00",
63404=>X"00",
63405=>X"00",
63406=>X"00",
63407=>X"00",
63408=>X"00",
63409=>X"00",
63410=>X"00",
63411=>X"00",
63412=>X"00",
63413=>X"00",
63414=>X"00",
63415=>X"00",
63416=>X"00",
63417=>X"00",
63418=>X"00",
63419=>X"00",
63420=>X"00",
63421=>X"00",
63422=>X"00",
63423=>X"00",
63424=>X"00",
63425=>X"00",
63426=>X"00",
63427=>X"00",
63428=>X"00",
63429=>X"00",
63430=>X"00",
63431=>X"00",
63432=>X"00",
63433=>X"00",
63434=>X"00",
63435=>X"00",
63436=>X"00",
63437=>X"00",
63438=>X"00",
63439=>X"00",
63440=>X"00",
63441=>X"00",
63442=>X"00",
63443=>X"00",
63444=>X"00",
63445=>X"00",
63446=>X"00",
63447=>X"00",
63448=>X"00",
63449=>X"00",
63450=>X"00",
63451=>X"00",
63452=>X"00",
63453=>X"00",
63454=>X"00",
63455=>X"00",
63456=>X"00",
63457=>X"00",
63458=>X"00",
63459=>X"00",
63460=>X"00",
63461=>X"00",
63462=>X"00",
63463=>X"00",
63464=>X"00",
63465=>X"00",
63466=>X"00",
63467=>X"00",
63468=>X"00",
63469=>X"00",
63470=>X"00",
63471=>X"00",
63472=>X"00",
63473=>X"00",
63474=>X"00",
63475=>X"00",
63476=>X"00",
63477=>X"00",
63478=>X"00",
63479=>X"00",
63480=>X"00",
63481=>X"00",
63482=>X"00",
63483=>X"00",
63484=>X"00",
63485=>X"00",
63486=>X"00",
63487=>X"00",
63488=>X"00",
63489=>X"00",
63490=>X"00",
63491=>X"00",
63492=>X"00",
63493=>X"00",
63494=>X"00",
63495=>X"00",
63496=>X"00",
63497=>X"00",
63498=>X"00",
63499=>X"00",
63500=>X"00",
63501=>X"00",
63502=>X"00",
63503=>X"00",
63504=>X"00",
63505=>X"00",
63506=>X"00",
63507=>X"00",
63508=>X"00",
63509=>X"00",
63510=>X"00",
63511=>X"00",
63512=>X"00",
63513=>X"00",
63514=>X"00",
63515=>X"00",
63516=>X"00",
63517=>X"00",
63518=>X"00",
63519=>X"00",
63520=>X"00",
63521=>X"00",
63522=>X"00",
63523=>X"00",
63524=>X"00",
63525=>X"00",
63526=>X"00",
63527=>X"00",
63528=>X"00",
63529=>X"00",
63530=>X"00",
63531=>X"00",
63532=>X"00",
63533=>X"00",
63534=>X"00",
63535=>X"00",
63536=>X"00",
63537=>X"00",
63538=>X"00",
63539=>X"00",
63540=>X"00",
63541=>X"00",
63542=>X"00",
63543=>X"00",
63544=>X"00",
63545=>X"00",
63546=>X"00",
63547=>X"00",
63548=>X"00",
63549=>X"00",
63550=>X"00",
63551=>X"00",
63552=>X"00",
63553=>X"00",
63554=>X"00",
63555=>X"00",
63556=>X"00",
63557=>X"00",
63558=>X"00",
63559=>X"00",
63560=>X"00",
63561=>X"00",
63562=>X"00",
63563=>X"00",
63564=>X"00",
63565=>X"00",
63566=>X"00",
63567=>X"00",
63568=>X"00",
63569=>X"00",
63570=>X"00",
63571=>X"00",
63572=>X"00",
63573=>X"00",
63574=>X"00",
63575=>X"00",
63576=>X"00",
63577=>X"00",
63578=>X"00",
63579=>X"00",
63580=>X"00",
63581=>X"00",
63582=>X"00",
63583=>X"00",
63584=>X"00",
63585=>X"00",
63586=>X"00",
63587=>X"00",
63588=>X"00",
63589=>X"00",
63590=>X"00",
63591=>X"00",
63592=>X"00",
63593=>X"00",
63594=>X"00",
63595=>X"00",
63596=>X"00",
63597=>X"00",
63598=>X"00",
63599=>X"00",
63600=>X"00",
63601=>X"00",
63602=>X"00",
63603=>X"00",
63604=>X"00",
63605=>X"00",
63606=>X"00",
63607=>X"00",
63608=>X"00",
63609=>X"00",
63610=>X"00",
63611=>X"00",
63612=>X"00",
63613=>X"00",
63614=>X"00",
63615=>X"00",
63616=>X"00",
63617=>X"00",
63618=>X"00",
63619=>X"00",
63620=>X"00",
63621=>X"00",
63622=>X"00",
63623=>X"00",
63624=>X"00",
63625=>X"00",
63626=>X"00",
63627=>X"00",
63628=>X"00",
63629=>X"00",
63630=>X"00",
63631=>X"00",
63632=>X"00",
63633=>X"00",
63634=>X"00",
63635=>X"00",
63636=>X"00",
63637=>X"00",
63638=>X"00",
63639=>X"00",
63640=>X"00",
63641=>X"00",
63642=>X"00",
63643=>X"00",
63644=>X"00",
63645=>X"00",
63646=>X"00",
63647=>X"00",
63648=>X"00",
63649=>X"00",
63650=>X"00",
63651=>X"00",
63652=>X"00",
63653=>X"00",
63654=>X"00",
63655=>X"00",
63656=>X"00",
63657=>X"00",
63658=>X"00",
63659=>X"00",
63660=>X"00",
63661=>X"00",
63662=>X"00",
63663=>X"00",
63664=>X"00",
63665=>X"00",
63666=>X"00",
63667=>X"00",
63668=>X"00",
63669=>X"00",
63670=>X"00",
63671=>X"00",
63672=>X"00",
63673=>X"00",
63674=>X"00",
63675=>X"00",
63676=>X"00",
63677=>X"00",
63678=>X"00",
63679=>X"00",
63680=>X"00",
63681=>X"00",
63682=>X"00",
63683=>X"00",
63684=>X"00",
63685=>X"00",
63686=>X"00",
63687=>X"00",
63688=>X"00",
63689=>X"00",
63690=>X"00",
63691=>X"00",
63692=>X"00",
63693=>X"00",
63694=>X"00",
63695=>X"00",
63696=>X"00",
63697=>X"00",
63698=>X"00",
63699=>X"00",
63700=>X"00",
63701=>X"00",
63702=>X"00",
63703=>X"00",
63704=>X"00",
63705=>X"00",
63706=>X"00",
63707=>X"00",
63708=>X"00",
63709=>X"00",
63710=>X"00",
63711=>X"00",
63712=>X"00",
63713=>X"00",
63714=>X"00",
63715=>X"00",
63716=>X"00",
63717=>X"00",
63718=>X"00",
63719=>X"00",
63720=>X"00",
63721=>X"00",
63722=>X"00",
63723=>X"00",
63724=>X"00",
63725=>X"00",
63726=>X"00",
63727=>X"00",
63728=>X"00",
63729=>X"00",
63730=>X"00",
63731=>X"00",
63732=>X"00",
63733=>X"00",
63734=>X"00",
63735=>X"00",
63736=>X"00",
63737=>X"00",
63738=>X"00",
63739=>X"00",
63740=>X"00",
63741=>X"00",
63742=>X"00",
63743=>X"00",
63744=>X"00",
63745=>X"00",
63746=>X"00",
63747=>X"00",
63748=>X"00",
63749=>X"00",
63750=>X"00",
63751=>X"00",
63752=>X"00",
63753=>X"00",
63754=>X"00",
63755=>X"00",
63756=>X"00",
63757=>X"00",
63758=>X"00",
63759=>X"00",
63760=>X"00",
63761=>X"00",
63762=>X"00",
63763=>X"00",
63764=>X"00",
63765=>X"00",
63766=>X"00",
63767=>X"00",
63768=>X"00",
63769=>X"00",
63770=>X"00",
63771=>X"00",
63772=>X"00",
63773=>X"00",
63774=>X"00",
63775=>X"00",
63776=>X"00",
63777=>X"00",
63778=>X"00",
63779=>X"00",
63780=>X"00",
63781=>X"00",
63782=>X"00",
63783=>X"00",
63784=>X"00",
63785=>X"00",
63786=>X"00",
63787=>X"00",
63788=>X"00",
63789=>X"00",
63790=>X"00",
63791=>X"00",
63792=>X"00",
63793=>X"00",
63794=>X"00",
63795=>X"00",
63796=>X"00",
63797=>X"00",
63798=>X"00",
63799=>X"00",
63800=>X"00",
63801=>X"00",
63802=>X"00",
63803=>X"00",
63804=>X"00",
63805=>X"00",
63806=>X"00",
63807=>X"00",
63808=>X"00",
63809=>X"00",
63810=>X"00",
63811=>X"00",
63812=>X"00",
63813=>X"00",
63814=>X"00",
63815=>X"00",
63816=>X"00",
63817=>X"00",
63818=>X"00",
63819=>X"00",
63820=>X"00",
63821=>X"00",
63822=>X"00",
63823=>X"00",
63824=>X"00",
63825=>X"00",
63826=>X"00",
63827=>X"00",
63828=>X"00",
63829=>X"00",
63830=>X"00",
63831=>X"00",
63832=>X"00",
63833=>X"00",
63834=>X"00",
63835=>X"00",
63836=>X"00",
63837=>X"00",
63838=>X"00",
63839=>X"00",
63840=>X"00",
63841=>X"00",
63842=>X"00",
63843=>X"00",
63844=>X"00",
63845=>X"00",
63846=>X"00",
63847=>X"00",
63848=>X"00",
63849=>X"00",
63850=>X"00",
63851=>X"00",
63852=>X"00",
63853=>X"00",
63854=>X"00",
63855=>X"00",
63856=>X"00",
63857=>X"00",
63858=>X"00",
63859=>X"00",
63860=>X"00",
63861=>X"00",
63862=>X"00",
63863=>X"00",
63864=>X"00",
63865=>X"00",
63866=>X"00",
63867=>X"00",
63868=>X"00",
63869=>X"00",
63870=>X"00",
63871=>X"00",
63872=>X"00",
63873=>X"00",
63874=>X"00",
63875=>X"00",
63876=>X"00",
63877=>X"00",
63878=>X"00",
63879=>X"00",
63880=>X"00",
63881=>X"00",
63882=>X"00",
63883=>X"00",
63884=>X"00",
63885=>X"00",
63886=>X"00",
63887=>X"00",
63888=>X"00",
63889=>X"00",
63890=>X"00",
63891=>X"00",
63892=>X"00",
63893=>X"00",
63894=>X"00",
63895=>X"00",
63896=>X"00",
63897=>X"00",
63898=>X"00",
63899=>X"00",
63900=>X"00",
63901=>X"00",
63902=>X"00",
63903=>X"00",
63904=>X"00",
63905=>X"00",
63906=>X"00",
63907=>X"00",
63908=>X"00",
63909=>X"00",
63910=>X"00",
63911=>X"00",
63912=>X"00",
63913=>X"00",
63914=>X"00",
63915=>X"00",
63916=>X"00",
63917=>X"00",
63918=>X"00",
63919=>X"00",
63920=>X"00",
63921=>X"00",
63922=>X"00",
63923=>X"00",
63924=>X"00",
63925=>X"00",
63926=>X"00",
63927=>X"00",
63928=>X"00",
63929=>X"00",
63930=>X"00",
63931=>X"00",
63932=>X"00",
63933=>X"00",
63934=>X"00",
63935=>X"00",
63936=>X"00",
63937=>X"00",
63938=>X"00",
63939=>X"00",
63940=>X"00",
63941=>X"00",
63942=>X"00",
63943=>X"00",
63944=>X"00",
63945=>X"00",
63946=>X"00",
63947=>X"00",
63948=>X"00",
63949=>X"00",
63950=>X"00",
63951=>X"00",
63952=>X"00",
63953=>X"00",
63954=>X"00",
63955=>X"00",
63956=>X"00",
63957=>X"00",
63958=>X"00",
63959=>X"00",
63960=>X"00",
63961=>X"00",
63962=>X"00",
63963=>X"00",
63964=>X"00",
63965=>X"00",
63966=>X"00",
63967=>X"00",
63968=>X"00",
63969=>X"00",
63970=>X"00",
63971=>X"00",
63972=>X"00",
63973=>X"00",
63974=>X"00",
63975=>X"00",
63976=>X"00",
63977=>X"00",
63978=>X"00",
63979=>X"00",
63980=>X"00",
63981=>X"00",
63982=>X"00",
63983=>X"00",
63984=>X"00",
63985=>X"00",
63986=>X"00",
63987=>X"00",
63988=>X"00",
63989=>X"00",
63990=>X"00",
63991=>X"00",
63992=>X"00",
63993=>X"00",
63994=>X"00",
63995=>X"00",
63996=>X"00",
63997=>X"00",
63998=>X"00",
63999=>X"00",
64000=>X"00",
64001=>X"00",
64002=>X"00",
64003=>X"00",
64004=>X"00",
64005=>X"00",
64006=>X"00",
64007=>X"00",
64008=>X"00",
64009=>X"00",
64010=>X"00",
64011=>X"00",
64012=>X"00",
64013=>X"00",
64014=>X"00",
64015=>X"00",
64016=>X"00",
64017=>X"00",
64018=>X"00",
64019=>X"00",
64020=>X"00",
64021=>X"00",
64022=>X"00",
64023=>X"00",
64024=>X"00",
64025=>X"00",
64026=>X"00",
64027=>X"00",
64028=>X"00",
64029=>X"00",
64030=>X"00",
64031=>X"00",
64032=>X"00",
64033=>X"00",
64034=>X"00",
64035=>X"00",
64036=>X"00",
64037=>X"00",
64038=>X"00",
64039=>X"00",
64040=>X"00",
64041=>X"00",
64042=>X"00",
64043=>X"00",
64044=>X"00",
64045=>X"00",
64046=>X"00",
64047=>X"00",
64048=>X"00",
64049=>X"00",
64050=>X"00",
64051=>X"00",
64052=>X"00",
64053=>X"00",
64054=>X"00",
64055=>X"00",
64056=>X"00",
64057=>X"00",
64058=>X"00",
64059=>X"00",
64060=>X"00",
64061=>X"00",
64062=>X"00",
64063=>X"00",
64064=>X"00",
64065=>X"00",
64066=>X"00",
64067=>X"00",
64068=>X"00",
64069=>X"00",
64070=>X"00",
64071=>X"00",
64072=>X"00",
64073=>X"00",
64074=>X"00",
64075=>X"00",
64076=>X"00",
64077=>X"00",
64078=>X"00",
64079=>X"00",
64080=>X"00",
64081=>X"00",
64082=>X"00",
64083=>X"00",
64084=>X"00",
64085=>X"00",
64086=>X"00",
64087=>X"00",
64088=>X"00",
64089=>X"00",
64090=>X"00",
64091=>X"00",
64092=>X"00",
64093=>X"00",
64094=>X"00",
64095=>X"00",
64096=>X"00",
64097=>X"00",
64098=>X"00",
64099=>X"00",
64100=>X"00",
64101=>X"00",
64102=>X"00",
64103=>X"00",
64104=>X"00",
64105=>X"00",
64106=>X"00",
64107=>X"00",
64108=>X"00",
64109=>X"00",
64110=>X"00",
64111=>X"00",
64112=>X"00",
64113=>X"00",
64114=>X"00",
64115=>X"00",
64116=>X"00",
64117=>X"00",
64118=>X"00",
64119=>X"00",
64120=>X"00",
64121=>X"00",
64122=>X"00",
64123=>X"00",
64124=>X"00",
64125=>X"00",
64126=>X"00",
64127=>X"00",
64128=>X"00",
64129=>X"00",
64130=>X"00",
64131=>X"00",
64132=>X"00",
64133=>X"00",
64134=>X"00",
64135=>X"00",
64136=>X"00",
64137=>X"00",
64138=>X"00",
64139=>X"00",
64140=>X"00",
64141=>X"00",
64142=>X"00",
64143=>X"00",
64144=>X"00",
64145=>X"00",
64146=>X"00",
64147=>X"00",
64148=>X"00",
64149=>X"00",
64150=>X"00",
64151=>X"00",
64152=>X"00",
64153=>X"00",
64154=>X"00",
64155=>X"00",
64156=>X"00",
64157=>X"00",
64158=>X"00",
64159=>X"00",
64160=>X"00",
64161=>X"00",
64162=>X"00",
64163=>X"00",
64164=>X"00",
64165=>X"00",
64166=>X"00",
64167=>X"00",
64168=>X"00",
64169=>X"00",
64170=>X"00",
64171=>X"00",
64172=>X"00",
64173=>X"00",
64174=>X"00",
64175=>X"00",
64176=>X"00",
64177=>X"00",
64178=>X"00",
64179=>X"00",
64180=>X"00",
64181=>X"00",
64182=>X"00",
64183=>X"00",
64184=>X"00",
64185=>X"00",
64186=>X"00",
64187=>X"00",
64188=>X"00",
64189=>X"00",
64190=>X"00",
64191=>X"00",
64192=>X"00",
64193=>X"00",
64194=>X"00",
64195=>X"00",
64196=>X"00",
64197=>X"00",
64198=>X"00",
64199=>X"00",
64200=>X"00",
64201=>X"00",
64202=>X"00",
64203=>X"00",
64204=>X"00",
64205=>X"00",
64206=>X"00",
64207=>X"00",
64208=>X"00",
64209=>X"00",
64210=>X"00",
64211=>X"00",
64212=>X"00",
64213=>X"00",
64214=>X"00",
64215=>X"00",
64216=>X"00",
64217=>X"00",
64218=>X"00",
64219=>X"00",
64220=>X"00",
64221=>X"00",
64222=>X"00",
64223=>X"00",
64224=>X"00",
64225=>X"00",
64226=>X"00",
64227=>X"00",
64228=>X"00",
64229=>X"00",
64230=>X"00",
64231=>X"00",
64232=>X"00",
64233=>X"00",
64234=>X"00",
64235=>X"00",
64236=>X"00",
64237=>X"00",
64238=>X"00",
64239=>X"00",
64240=>X"00",
64241=>X"00",
64242=>X"00",
64243=>X"00",
64244=>X"00",
64245=>X"00",
64246=>X"00",
64247=>X"00",
64248=>X"00",
64249=>X"00",
64250=>X"00",
64251=>X"00",
64252=>X"00",
64253=>X"00",
64254=>X"00",
64255=>X"00",
64256=>X"00",
64257=>X"00",
64258=>X"00",
64259=>X"00",
64260=>X"00",
64261=>X"00",
64262=>X"00",
64263=>X"00",
64264=>X"00",
64265=>X"00",
64266=>X"00",
64267=>X"00",
64268=>X"00",
64269=>X"00",
64270=>X"00",
64271=>X"00",
64272=>X"00",
64273=>X"00",
64274=>X"00",
64275=>X"00",
64276=>X"00",
64277=>X"00",
64278=>X"00",
64279=>X"00",
64280=>X"00",
64281=>X"00",
64282=>X"00",
64283=>X"00",
64284=>X"00",
64285=>X"00",
64286=>X"00",
64287=>X"00",
64288=>X"00",
64289=>X"00",
64290=>X"00",
64291=>X"00",
64292=>X"00",
64293=>X"00",
64294=>X"00",
64295=>X"00",
64296=>X"00",
64297=>X"00",
64298=>X"00",
64299=>X"00",
64300=>X"00",
64301=>X"00",
64302=>X"00",
64303=>X"00",
64304=>X"00",
64305=>X"00",
64306=>X"00",
64307=>X"00",
64308=>X"00",
64309=>X"00",
64310=>X"00",
64311=>X"00",
64312=>X"00",
64313=>X"00",
64314=>X"00",
64315=>X"00",
64316=>X"00",
64317=>X"00",
64318=>X"00",
64319=>X"00",
64320=>X"00",
64321=>X"00",
64322=>X"00",
64323=>X"00",
64324=>X"00",
64325=>X"00",
64326=>X"00",
64327=>X"00",
64328=>X"00",
64329=>X"00",
64330=>X"00",
64331=>X"00",
64332=>X"00",
64333=>X"00",
64334=>X"00",
64335=>X"00",
64336=>X"00",
64337=>X"00",
64338=>X"00",
64339=>X"00",
64340=>X"00",
64341=>X"00",
64342=>X"00",
64343=>X"00",
64344=>X"00",
64345=>X"00",
64346=>X"00",
64347=>X"00",
64348=>X"00",
64349=>X"00",
64350=>X"00",
64351=>X"00",
64352=>X"00",
64353=>X"00",
64354=>X"00",
64355=>X"00",
64356=>X"00",
64357=>X"00",
64358=>X"00",
64359=>X"00",
64360=>X"00",
64361=>X"00",
64362=>X"00",
64363=>X"00",
64364=>X"00",
64365=>X"00",
64366=>X"00",
64367=>X"00",
64368=>X"00",
64369=>X"00",
64370=>X"00",
64371=>X"00",
64372=>X"00",
64373=>X"00",
64374=>X"00",
64375=>X"00",
64376=>X"00",
64377=>X"00",
64378=>X"00",
64379=>X"00",
64380=>X"00",
64381=>X"00",
64382=>X"00",
64383=>X"00",
64384=>X"00",
64385=>X"00",
64386=>X"00",
64387=>X"00",
64388=>X"00",
64389=>X"00",
64390=>X"00",
64391=>X"00",
64392=>X"00",
64393=>X"00",
64394=>X"00",
64395=>X"00",
64396=>X"00",
64397=>X"00",
64398=>X"00",
64399=>X"00",
64400=>X"00",
64401=>X"00",
64402=>X"00",
64403=>X"00",
64404=>X"00",
64405=>X"00",
64406=>X"00",
64407=>X"00",
64408=>X"00",
64409=>X"00",
64410=>X"00",
64411=>X"00",
64412=>X"00",
64413=>X"00",
64414=>X"00",
64415=>X"00",
64416=>X"00",
64417=>X"00",
64418=>X"00",
64419=>X"00",
64420=>X"00",
64421=>X"00",
64422=>X"00",
64423=>X"00",
64424=>X"00",
64425=>X"00",
64426=>X"00",
64427=>X"00",
64428=>X"00",
64429=>X"00",
64430=>X"00",
64431=>X"00",
64432=>X"00",
64433=>X"00",
64434=>X"00",
64435=>X"00",
64436=>X"00",
64437=>X"00",
64438=>X"00",
64439=>X"00",
64440=>X"00",
64441=>X"00",
64442=>X"00",
64443=>X"00",
64444=>X"00",
64445=>X"00",
64446=>X"00",
64447=>X"00",
64448=>X"00",
64449=>X"00",
64450=>X"00",
64451=>X"00",
64452=>X"00",
64453=>X"00",
64454=>X"00",
64455=>X"00",
64456=>X"00",
64457=>X"00",
64458=>X"00",
64459=>X"00",
64460=>X"00",
64461=>X"00",
64462=>X"00",
64463=>X"00",
64464=>X"00",
64465=>X"00",
64466=>X"00",
64467=>X"00",
64468=>X"00",
64469=>X"00",
64470=>X"00",
64471=>X"00",
64472=>X"00",
64473=>X"00",
64474=>X"00",
64475=>X"00",
64476=>X"00",
64477=>X"00",
64478=>X"00",
64479=>X"00",
64480=>X"00",
64481=>X"00",
64482=>X"00",
64483=>X"00",
64484=>X"00",
64485=>X"00",
64486=>X"00",
64487=>X"00",
64488=>X"00",
64489=>X"00",
64490=>X"00",
64491=>X"00",
64492=>X"00",
64493=>X"00",
64494=>X"00",
64495=>X"00",
64496=>X"00",
64497=>X"00",
64498=>X"00",
64499=>X"00",
64500=>X"00",
64501=>X"00",
64502=>X"00",
64503=>X"00",
64504=>X"00",
64505=>X"00",
64506=>X"00",
64507=>X"00",
64508=>X"00",
64509=>X"00",
64510=>X"00",
64511=>X"00",
64512=>X"00",
64513=>X"00",
64514=>X"00",
64515=>X"00",
64516=>X"00",
64517=>X"00",
64518=>X"00",
64519=>X"00",
64520=>X"00",
64521=>X"00",
64522=>X"00",
64523=>X"00",
64524=>X"00",
64525=>X"00",
64526=>X"00",
64527=>X"00",
64528=>X"00",
64529=>X"00",
64530=>X"00",
64531=>X"00",
64532=>X"00",
64533=>X"00",
64534=>X"00",
64535=>X"00",
64536=>X"00",
64537=>X"00",
64538=>X"00",
64539=>X"00",
64540=>X"00",
64541=>X"00",
64542=>X"00",
64543=>X"00",
64544=>X"00",
64545=>X"00",
64546=>X"00",
64547=>X"00",
64548=>X"00",
64549=>X"00",
64550=>X"00",
64551=>X"00",
64552=>X"00",
64553=>X"00",
64554=>X"00",
64555=>X"00",
64556=>X"00",
64557=>X"00",
64558=>X"00",
64559=>X"00",
64560=>X"00",
64561=>X"00",
64562=>X"00",
64563=>X"00",
64564=>X"00",
64565=>X"00",
64566=>X"00",
64567=>X"00",
64568=>X"00",
64569=>X"00",
64570=>X"00",
64571=>X"00",
64572=>X"00",
64573=>X"00",
64574=>X"00",
64575=>X"00",
64576=>X"00",
64577=>X"00",
64578=>X"00",
64579=>X"00",
64580=>X"00",
64581=>X"00",
64582=>X"00",
64583=>X"00",
64584=>X"00",
64585=>X"00",
64586=>X"00",
64587=>X"00",
64588=>X"00",
64589=>X"00",
64590=>X"00",
64591=>X"00",
64592=>X"00",
64593=>X"00",
64594=>X"00",
64595=>X"00",
64596=>X"00",
64597=>X"00",
64598=>X"00",
64599=>X"00",
64600=>X"00",
64601=>X"00",
64602=>X"00",
64603=>X"00",
64604=>X"00",
64605=>X"00",
64606=>X"00",
64607=>X"00",
64608=>X"00",
64609=>X"00",
64610=>X"00",
64611=>X"00",
64612=>X"00",
64613=>X"00",
64614=>X"00",
64615=>X"00",
64616=>X"00",
64617=>X"00",
64618=>X"00",
64619=>X"00",
64620=>X"00",
64621=>X"00",
64622=>X"00",
64623=>X"00",
64624=>X"00",
64625=>X"00",
64626=>X"00",
64627=>X"00",
64628=>X"00",
64629=>X"00",
64630=>X"00",
64631=>X"00",
64632=>X"00",
64633=>X"00",
64634=>X"00",
64635=>X"00",
64636=>X"00",
64637=>X"00",
64638=>X"00",
64639=>X"00",
64640=>X"00",
64641=>X"00",
64642=>X"00",
64643=>X"00",
64644=>X"00",
64645=>X"00",
64646=>X"00",
64647=>X"00",
64648=>X"00",
64649=>X"00",
64650=>X"00",
64651=>X"00",
64652=>X"00",
64653=>X"00",
64654=>X"00",
64655=>X"00",
64656=>X"00",
64657=>X"00",
64658=>X"00",
64659=>X"00",
64660=>X"00",
64661=>X"00",
64662=>X"00",
64663=>X"00",
64664=>X"00",
64665=>X"00",
64666=>X"00",
64667=>X"00",
64668=>X"00",
64669=>X"00",
64670=>X"00",
64671=>X"00",
64672=>X"00",
64673=>X"00",
64674=>X"00",
64675=>X"00",
64676=>X"00",
64677=>X"00",
64678=>X"00",
64679=>X"00",
64680=>X"00",
64681=>X"00",
64682=>X"00",
64683=>X"00",
64684=>X"00",
64685=>X"00",
64686=>X"00",
64687=>X"00",
64688=>X"00",
64689=>X"00",
64690=>X"00",
64691=>X"00",
64692=>X"00",
64693=>X"00",
64694=>X"00",
64695=>X"00",
64696=>X"00",
64697=>X"00",
64698=>X"00",
64699=>X"00",
64700=>X"00",
64701=>X"00",
64702=>X"00",
64703=>X"00",
64704=>X"00",
64705=>X"00",
64706=>X"00",
64707=>X"00",
64708=>X"00",
64709=>X"00",
64710=>X"00",
64711=>X"00",
64712=>X"00",
64713=>X"00",
64714=>X"00",
64715=>X"00",
64716=>X"00",
64717=>X"00",
64718=>X"00",
64719=>X"00",
64720=>X"00",
64721=>X"00",
64722=>X"00",
64723=>X"00",
64724=>X"00",
64725=>X"00",
64726=>X"00",
64727=>X"00",
64728=>X"00",
64729=>X"00",
64730=>X"00",
64731=>X"00",
64732=>X"00",
64733=>X"00",
64734=>X"00",
64735=>X"00",
64736=>X"00",
64737=>X"00",
64738=>X"00",
64739=>X"00",
64740=>X"00",
64741=>X"00",
64742=>X"00",
64743=>X"00",
64744=>X"00",
64745=>X"00",
64746=>X"00",
64747=>X"00",
64748=>X"00",
64749=>X"00",
64750=>X"00",
64751=>X"00",
64752=>X"00",
64753=>X"00",
64754=>X"00",
64755=>X"00",
64756=>X"00",
64757=>X"00",
64758=>X"00",
64759=>X"00",
64760=>X"00",
64761=>X"00",
64762=>X"00",
64763=>X"00",
64764=>X"00",
64765=>X"00",
64766=>X"00",
64767=>X"00",
64768=>X"00",
64769=>X"00",
64770=>X"00",
64771=>X"00",
64772=>X"00",
64773=>X"00",
64774=>X"00",
64775=>X"00",
64776=>X"00",
64777=>X"00",
64778=>X"00",
64779=>X"00",
64780=>X"00",
64781=>X"00",
64782=>X"00",
64783=>X"00",
64784=>X"00",
64785=>X"00",
64786=>X"00",
64787=>X"00",
64788=>X"00",
64789=>X"00",
64790=>X"00",
64791=>X"00",
64792=>X"00",
64793=>X"00",
64794=>X"00",
64795=>X"00",
64796=>X"00",
64797=>X"00",
64798=>X"00",
64799=>X"00",
64800=>X"00",
64801=>X"00",
64802=>X"00",
64803=>X"00",
64804=>X"00",
64805=>X"00",
64806=>X"00",
64807=>X"00",
64808=>X"00",
64809=>X"00",
64810=>X"00",
64811=>X"00",
64812=>X"00",
64813=>X"00",
64814=>X"00",
64815=>X"00",
64816=>X"00",
64817=>X"00",
64818=>X"00",
64819=>X"00",
64820=>X"00",
64821=>X"00",
64822=>X"00",
64823=>X"00",
64824=>X"00",
64825=>X"00",
64826=>X"00",
64827=>X"00",
64828=>X"00",
64829=>X"00",
64830=>X"00",
64831=>X"00",
64832=>X"00",
64833=>X"00",
64834=>X"00",
64835=>X"00",
64836=>X"00",
64837=>X"00",
64838=>X"00",
64839=>X"00",
64840=>X"00",
64841=>X"00",
64842=>X"00",
64843=>X"00",
64844=>X"00",
64845=>X"00",
64846=>X"00",
64847=>X"00",
64848=>X"00",
64849=>X"00",
64850=>X"00",
64851=>X"00",
64852=>X"00",
64853=>X"00",
64854=>X"00",
64855=>X"00",
64856=>X"00",
64857=>X"00",
64858=>X"00",
64859=>X"00",
64860=>X"00",
64861=>X"00",
64862=>X"00",
64863=>X"00",
64864=>X"00",
64865=>X"00",
64866=>X"00",
64867=>X"00",
64868=>X"00",
64869=>X"00",
64870=>X"00",
64871=>X"00",
64872=>X"00",
64873=>X"00",
64874=>X"00",
64875=>X"00",
64876=>X"00",
64877=>X"00",
64878=>X"00",
64879=>X"00",
64880=>X"00",
64881=>X"00",
64882=>X"00",
64883=>X"00",
64884=>X"00",
64885=>X"00",
64886=>X"00",
64887=>X"00",
64888=>X"00",
64889=>X"00",
64890=>X"00",
64891=>X"00",
64892=>X"00",
64893=>X"00",
64894=>X"00",
64895=>X"00",
64896=>X"00",
64897=>X"00",
64898=>X"00",
64899=>X"00",
64900=>X"00",
64901=>X"00",
64902=>X"00",
64903=>X"00",
64904=>X"00",
64905=>X"00",
64906=>X"00",
64907=>X"00",
64908=>X"00",
64909=>X"00",
64910=>X"00",
64911=>X"00",
64912=>X"00",
64913=>X"00",
64914=>X"00",
64915=>X"00",
64916=>X"00",
64917=>X"00",
64918=>X"00",
64919=>X"00",
64920=>X"00",
64921=>X"00",
64922=>X"00",
64923=>X"00",
64924=>X"00",
64925=>X"00",
64926=>X"00",
64927=>X"00",
64928=>X"00",
64929=>X"00",
64930=>X"00",
64931=>X"00",
64932=>X"00",
64933=>X"00",
64934=>X"00",
64935=>X"00",
64936=>X"00",
64937=>X"00",
64938=>X"00",
64939=>X"00",
64940=>X"00",
64941=>X"00",
64942=>X"00",
64943=>X"00",
64944=>X"00",
64945=>X"00",
64946=>X"00",
64947=>X"00",
64948=>X"00",
64949=>X"00",
64950=>X"00",
64951=>X"00",
64952=>X"00",
64953=>X"00",
64954=>X"00",
64955=>X"00",
64956=>X"00",
64957=>X"00",
64958=>X"00",
64959=>X"00",
64960=>X"00",
64961=>X"00",
64962=>X"00",
64963=>X"00",
64964=>X"00",
64965=>X"00",
64966=>X"00",
64967=>X"00",
64968=>X"00",
64969=>X"00",
64970=>X"00",
64971=>X"00",
64972=>X"00",
64973=>X"00",
64974=>X"00",
64975=>X"00",
64976=>X"00",
64977=>X"00",
64978=>X"00",
64979=>X"00",
64980=>X"00",
64981=>X"00",
64982=>X"00",
64983=>X"00",
64984=>X"00",
64985=>X"00",
64986=>X"00",
64987=>X"00",
64988=>X"00",
64989=>X"00",
64990=>X"00",
64991=>X"00",
64992=>X"00",
64993=>X"00",
64994=>X"00",
64995=>X"00",
64996=>X"00",
64997=>X"00",
64998=>X"00",
64999=>X"00",
65000=>X"00",
65001=>X"00",
65002=>X"00",
65003=>X"00",
65004=>X"00",
65005=>X"00",
65006=>X"00",
65007=>X"00",
65008=>X"00",
65009=>X"00",
65010=>X"00",
65011=>X"00",
65012=>X"00",
65013=>X"00",
65014=>X"00",
65015=>X"00",
65016=>X"00",
65017=>X"00",
65018=>X"00",
65019=>X"00",
65020=>X"00",
65021=>X"00",
65022=>X"00",
65023=>X"00",
65024=>X"00",
65025=>X"00",
65026=>X"00",
65027=>X"00",
65028=>X"00",
65029=>X"00",
65030=>X"00",
65031=>X"00",
65032=>X"00",
65033=>X"00",
65034=>X"00",
65035=>X"00",
65036=>X"00",
65037=>X"00",
65038=>X"00",
65039=>X"00",
65040=>X"00",
65041=>X"00",
65042=>X"00",
65043=>X"00",
65044=>X"00",
65045=>X"00",
65046=>X"00",
65047=>X"00",
65048=>X"00",
65049=>X"00",
65050=>X"00",
65051=>X"00",
65052=>X"00",
65053=>X"00",
65054=>X"00",
65055=>X"00",
65056=>X"00",
65057=>X"00",
65058=>X"00",
65059=>X"00",
65060=>X"00",
65061=>X"00",
65062=>X"00",
65063=>X"00",
65064=>X"00",
65065=>X"00",
65066=>X"00",
65067=>X"00",
65068=>X"00",
65069=>X"00",
65070=>X"00",
65071=>X"00",
65072=>X"00",
65073=>X"00",
65074=>X"00",
65075=>X"00",
65076=>X"00",
65077=>X"00",
65078=>X"00",
65079=>X"00",
65080=>X"00",
65081=>X"00",
65082=>X"00",
65083=>X"00",
65084=>X"00",
65085=>X"00",
65086=>X"00",
65087=>X"00",
65088=>X"00",
65089=>X"00",
65090=>X"00",
65091=>X"00",
65092=>X"00",
65093=>X"00",
65094=>X"00",
65095=>X"00",
65096=>X"00",
65097=>X"00",
65098=>X"00",
65099=>X"00",
65100=>X"00",
65101=>X"00",
65102=>X"00",
65103=>X"00",
65104=>X"00",
65105=>X"00",
65106=>X"00",
65107=>X"00",
65108=>X"00",
65109=>X"00",
65110=>X"00",
65111=>X"00",
65112=>X"00",
65113=>X"00",
65114=>X"00",
65115=>X"00",
65116=>X"00",
65117=>X"00",
65118=>X"00",
65119=>X"00",
65120=>X"00",
65121=>X"00",
65122=>X"00",
65123=>X"00",
65124=>X"00",
65125=>X"00",
65126=>X"00",
65127=>X"00",
65128=>X"00",
65129=>X"00",
65130=>X"00",
65131=>X"00",
65132=>X"00",
65133=>X"00",
65134=>X"00",
65135=>X"00",
65136=>X"00",
65137=>X"00",
65138=>X"00",
65139=>X"00",
65140=>X"00",
65141=>X"00",
65142=>X"00",
65143=>X"00",
65144=>X"00",
65145=>X"00",
65146=>X"00",
65147=>X"00",
65148=>X"00",
65149=>X"00",
65150=>X"00",
65151=>X"00",
65152=>X"00",
65153=>X"00",
65154=>X"00",
65155=>X"00",
65156=>X"00",
65157=>X"00",
65158=>X"00",
65159=>X"00",
65160=>X"00",
65161=>X"00",
65162=>X"00",
65163=>X"00",
65164=>X"00",
65165=>X"00",
65166=>X"00",
65167=>X"00",
65168=>X"00",
65169=>X"00",
65170=>X"00",
65171=>X"00",
65172=>X"00",
65173=>X"00",
65174=>X"00",
65175=>X"00",
65176=>X"00",
65177=>X"00",
65178=>X"00",
65179=>X"00",
65180=>X"00",
65181=>X"00",
65182=>X"00",
65183=>X"00",
65184=>X"00",
65185=>X"00",
65186=>X"00",
65187=>X"00",
65188=>X"00",
65189=>X"00",
65190=>X"00",
65191=>X"00",
65192=>X"00",
65193=>X"00",
65194=>X"00",
65195=>X"00",
65196=>X"00",
65197=>X"00",
65198=>X"00",
65199=>X"00",
65200=>X"00",
65201=>X"00",
65202=>X"00",
65203=>X"00",
65204=>X"00",
65205=>X"00",
65206=>X"00",
65207=>X"00",
65208=>X"00",
65209=>X"00",
65210=>X"00",
65211=>X"00",
65212=>X"00",
65213=>X"00",
65214=>X"00",
65215=>X"00",
65216=>X"00",
65217=>X"00",
65218=>X"00",
65219=>X"00",
65220=>X"00",
65221=>X"00",
65222=>X"00",
65223=>X"00",
65224=>X"00",
65225=>X"00",
65226=>X"00",
65227=>X"00",
65228=>X"00",
65229=>X"00",
65230=>X"00",
65231=>X"00",
65232=>X"00",
65233=>X"00",
65234=>X"00",
65235=>X"00",
65236=>X"00",
65237=>X"00",
65238=>X"00",
65239=>X"00",
65240=>X"00",
65241=>X"00",
65242=>X"00",
65243=>X"00",
65244=>X"00",
65245=>X"00",
65246=>X"00",
65247=>X"00",
65248=>X"00",
65249=>X"00",
65250=>X"00",
65251=>X"00",
65252=>X"00",
65253=>X"00",
65254=>X"00",
65255=>X"00",
65256=>X"00",
65257=>X"00",
65258=>X"00",
65259=>X"00",
65260=>X"00",
65261=>X"00",
65262=>X"00",
65263=>X"00",
65264=>X"00",
65265=>X"00",
65266=>X"00",
65267=>X"00",
65268=>X"00",
65269=>X"00",
65270=>X"00",
65271=>X"00",
65272=>X"00",
65273=>X"00",
65274=>X"00",
65275=>X"00",
65276=>X"00",
65277=>X"00",
65278=>X"00",
65279=>X"00",
65280=>X"00",
65281=>X"00",
65282=>X"00",
65283=>X"00",
65284=>X"00",
65285=>X"00",
65286=>X"00",
65287=>X"00",
65288=>X"00",
65289=>X"00",
65290=>X"00",
65291=>X"00",
65292=>X"00",
65293=>X"00",
65294=>X"00",
65295=>X"00",
65296=>X"00",
65297=>X"00",
65298=>X"00",
65299=>X"00",
65300=>X"00",
65301=>X"00",
65302=>X"00",
65303=>X"00",
65304=>X"00",
65305=>X"00",
65306=>X"00",
65307=>X"00",
65308=>X"00",
65309=>X"00",
65310=>X"00",
65311=>X"00",
65312=>X"00",
65313=>X"00",
65314=>X"00",
65315=>X"00",
65316=>X"00",
65317=>X"00",
65318=>X"00",
65319=>X"00",
65320=>X"00",
65321=>X"00",
65322=>X"00",
65323=>X"00",
65324=>X"00",
65325=>X"00",
65326=>X"00",
65327=>X"00",
65328=>X"00",
65329=>X"00",
65330=>X"00",
65331=>X"00",
65332=>X"00",
65333=>X"00",
65334=>X"00",
65335=>X"00",
65336=>X"00",
65337=>X"00",
65338=>X"00",
65339=>X"00",
65340=>X"00",
65341=>X"00",
65342=>X"00",
65343=>X"00",
65344=>X"00",
65345=>X"00",
65346=>X"00",
65347=>X"00",
65348=>X"00",
65349=>X"00",
65350=>X"00",
65351=>X"00",
65352=>X"00",
65353=>X"00",
65354=>X"00",
65355=>X"00",
65356=>X"00",
65357=>X"00",
65358=>X"00",
65359=>X"00",
65360=>X"00",
65361=>X"00",
65362=>X"00",
65363=>X"00",
65364=>X"00",
65365=>X"00",
65366=>X"00",
65367=>X"00",
65368=>X"00",
65369=>X"00",
65370=>X"00",
65371=>X"00",
65372=>X"00",
65373=>X"00",
65374=>X"00",
65375=>X"00",
65376=>X"00",
65377=>X"00",
65378=>X"00",
65379=>X"00",
65380=>X"00",
65381=>X"00",
65382=>X"00",
65383=>X"00",
65384=>X"00",
65385=>X"00",
65386=>X"00",
65387=>X"00",
65388=>X"00",
65389=>X"00",
65390=>X"00",
65391=>X"00",
65392=>X"00",
65393=>X"00",
65394=>X"00",
65395=>X"00",
65396=>X"00",
65397=>X"00",
65398=>X"00",
65399=>X"00",
65400=>X"00",
65401=>X"00",
65402=>X"00",
65403=>X"00",
65404=>X"00",
65405=>X"00",
65406=>X"00",
65407=>X"00",
65408=>X"00",
65409=>X"00",
65410=>X"00",
65411=>X"00",
65412=>X"00",
65413=>X"00",
65414=>X"00",
65415=>X"00",
65416=>X"00",
65417=>X"00",
65418=>X"00",
65419=>X"00",
65420=>X"00",
65421=>X"00",
65422=>X"00",
65423=>X"00",
65424=>X"00",
65425=>X"00",
65426=>X"00",
65427=>X"00",
65428=>X"00",
65429=>X"00",
65430=>X"00",
65431=>X"00",
65432=>X"00",
65433=>X"00",
65434=>X"00",
65435=>X"00",
65436=>X"00",
65437=>X"00",
65438=>X"00",
65439=>X"00",
65440=>X"00",
65441=>X"00",
65442=>X"00",
65443=>X"00",
65444=>X"00",
65445=>X"00",
65446=>X"00",
65447=>X"00",
65448=>X"00",
65449=>X"00",
65450=>X"00",
65451=>X"00",
65452=>X"00",
65453=>X"00",
65454=>X"00",
65455=>X"00",
65456=>X"00",
65457=>X"00",
65458=>X"00",
65459=>X"00",
65460=>X"00",
65461=>X"00",
65462=>X"00",
65463=>X"00",
65464=>X"00",
65465=>X"00",
65466=>X"00",
65467=>X"00",
65468=>X"00",
65469=>X"00",
65470=>X"00",
65471=>X"00",
65472=>X"00",
65473=>X"00",
65474=>X"00",
65475=>X"00",
65476=>X"00",
65477=>X"00",
65478=>X"00",
65479=>X"00",
65480=>X"00",
65481=>X"00",
65482=>X"00",
65483=>X"00",
65484=>X"00",
65485=>X"00",
65486=>X"00",
65487=>X"00",
65488=>X"00",
65489=>X"00",
65490=>X"00",
65491=>X"00",
65492=>X"00",
65493=>X"00",
65494=>X"00",
65495=>X"00",
65496=>X"00",
65497=>X"00",
65498=>X"00",
65499=>X"00",
65500=>X"00",
65501=>X"00",
65502=>X"00",
65503=>X"00",
65504=>X"00",
65505=>X"00",
65506=>X"00",
65507=>X"00",
65508=>X"00",
65509=>X"00",
65510=>X"00",
65511=>X"00",
65512=>X"00",
65513=>X"00",
65514=>X"00",
65515=>X"00",
65516=>X"00",
65517=>X"00",
65518=>X"00",
65519=>X"00",
65520=>X"00",
65521=>X"00",
65522=>X"00",
65523=>X"00",
65524=>X"00",
65525=>X"00",
65526=>X"00",
65527=>X"00",
65528=>X"00",
65529=>X"00",
65530=>X"00",
65531=>X"00",
65532=>X"00",
65533=>X"00",
65534=>X"00",
65535=>X"00",
     others => X"00");
attribute rom_block: string;
attribute rom_block of ROMINIT : constant is "ROM_CELL_XYZ01";
begin

process
begin
  wait until rising_edge(clk_25);

  if (reset='1') then
    h_count     <= "0000000000";
	v_count     <= "0000000000";
	new_frame   <= '0';
    frame_num   <= "0111110100";
  else
	
	new_frame  <= '0'; -- default
	if (h_count = "1100011111") then
	  h_count <= "0000000000";
	  if ( v_count = "1000001100" ) then
        v_count     <= "0000000000";
        new_frame   <= '0';                
      else
        v_count <= v_count + 1;
      end if; -- v_count
    else  
      h_count <= h_count + 1;
    end if; -- h_count
        
    if (new_frame = '1') then
      if (frame_num = "1111111111") then
        frame_num <= "0000000000";
      else
        frame_num <= frame_num + 1;
      end if;
    end if;
  end if; -- reset
end process;  
Leer:process(h_count, v_count)
variable direcciones: std_logic_vector(13 downto 0):="00000000000000";
variable valores_totales: std_logic_vector(7 downto 0);
begin
direcciones( 6 downto 0):=h_count(7 downto 1);
direcciones( 13 downto 7):=v_count(8 downto 2);
valores_totales := ROMINIT(TO_INTEGER(UNSIGNED(direcciones)));

 if ( h_count < "01100000" ) then
    hs_1 <= '1';  else
    hs_1 <= '0';  end if;

  if ( v_count <"000000010") then
    vs_1 <= '1';  else
    vs_1 <= '0';  end if;

  if ( h_count >= "0010010000") and
     ( h_count <  "1100010000" ) and
     ( v_count >= "0000100100" ) and
     ( v_count <  "1000000100" ) then
    de_1 <= '1'; else
    de_1 <= '0'; end if;
hs_out  <= hs_1;
vs_out  <= vs_1;
r_out   <= valores_totales(5 downto 4);
de_out  <= de_1;
g_out   <= valores_totales(3 downto  2);
b_out   <= valores_totales(1 downto  0);
end process;

end behave;